// Verilog netlist created by TD v4.4.433
// Fri May 10 11:03:38 2019

`timescale 1ns / 1ps
module ImgROM  // al_ip/ROM.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [14:0] addra;  // al_ip/ROM.v(18)
  input clka;  // al_ip/ROM.v(19)
  input rsta;  // al_ip/ROM.v(20)
  output [7:0] doa;  // al_ip/ROM.v(16)

  wire [0:1] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;

  reg_sr_as_w1 addra_pipe_b0 (
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[0]));
  reg_sr_as_w1 addra_pipe_b1 (
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .reset(rsta),
    .set(1'b0),
    .q(addra_piped[1]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFCD565FBD6555555555C77FC15DBA7DDF77FCF5555555555555555555D7E036),
    .INIT_01(256'hFF57F75E390FFFFFFFFF7F47A1FF73FD1D74FDDFFFFFFFF5FDFFDFFFF6CE2FBE),
    .INIT_02(256'hFF4F7D7DDD5FFFFFFFFD7F4535D18E1D9551575FFFFD7776D0D55EB43F6F3F41),
    .INIT_03(256'hFF6F5F5B7E5FFFFFFFFFEF6C05D6D15D956DEFF5FFF5F3B76BA0B1A641FD772F),
    .INIT_04(256'hFF4DE5F9C47FFFFFFFFF074ED547DF8D11CDFFF5FFD436497F3FDE5F57DD60F7),
    .INIT_05(256'hFF4D1FFC45DFFFFFD5F6174C9DE242EDD39DBFFFFFDBA7FD0433435FDFF71BFF),
    .INIT_06(256'hFF6D95DDE77FFFFFD5FDFD7A5D37F565D956FFFFFFDDFD3AB9DE35FFFDD5BFFF),
    .INIT_07(256'hFF4F71FEB7FFFFFFD5FF75B9755C78A9525D7FFFFFF775B35F8D7FFFFD60DFFF),
    .INIT_08(256'hFF57FFFF9FFFD5FFD55C1F125437FC2353D9FFFF75D9D9DF5A57FFFFFF77F618),
    .INIT_09(256'hFFD7D3FF4FFFFD7FD558FD2B5A4E3E4A7FFBFFFFFEFC7F5C157FD7FFFF5D6AC3),
    .INIT_0A(256'hFFC5EDDD67FFFC5FD5F1FD857D8DDD3DFFE7FFF56315D70D7FF557FFFD77C002),
    .INIT_0B(256'hFF615BDDDFFFD497D7FFFD194EFDAF167F77F7F75DF77A5FFFFD57FD7FDA0A55),
    .INIT_0C(256'hFFDB485E5FFFC5D97FF67D5B961FF7733D17F5D47FFEBD5555557FFFFFDE7FFF),
    .INIT_0D(256'hFFD759DDFD7F4EFE5F7E750DBDA5DF4E3D97F54DFFDE800002A355FFFFF7FFFF),
    .INIT_0E(256'hFFC57CDF59D7DB1D6D5F559DF9D829E33C75D657FFF55555555DCA555FFDFFFF),
    .INIT_0F(256'hFFD37D747717D451F9EF56EC60FFF5E8F65F797FFFFDFFFFFFFF55D857F758FF),
    .INIT_10(256'hCDCDD8767D4955D57FB356F4F41A22A2D957BFFC15FFFFFFFFFFFF55C955DE8F),
    .INIT_11(256'hD57054D47FD69597F57F76BDD4FC2FE0D15D70530C7FFFFFFFFFFFFFF7A5775B),
    .INIT_12(256'hBE5EDD167FFFC9ED7C997731E0C35173554BB1B159DF0A9FFFFFFFFFF5F495E5),
    .INIT_13(256'hAF2E77C5FFFFF72319057D71067A621AC5562F23C25602C7709FFFFFF020B5D4),
    .INIT_14(256'h6969DE7F9FFFFF7F4D35FCBF338D6B88799C98A726EEB0BFC5E69555755555F5),
    .INIT_15(256'hCBD47D7B9FFFDFDFD9FF56AE2D18A16D3F34DD6575DF60BFF4A0AF357FFD7FF5),
    .INIT_16(256'hF3DCB7AD77FFFD7C5F3F5E5D87FFDFF2B75D7FFD57DF3683FFFF72CFA77FFFFF),
    .INIT_17(256'hF79D97EEC7FFFFCC273F5D7E5FFFFFFD5FDDFFFFFFD5D2413FFFFF5A051D5FFF),
    .INIT_18(256'hFF555D0D47FFFC7227EF55321FFFFFFD555DFFFFFFF5774DD3FFFFD5D42CF5F7),
    .INIT_19(256'hFF5DF54597FFF73EF46F4D1E5D7FFFFD557FFFFFFFFFFC8F4FFFFFFFFFF37355),
    .INIT_1A(256'hFFAFFD5DD7FFDAC5D47FA5D15D7FFFFFF57FFFFFFFFD7DA530FFFFFFFFFD5EC5),
    .INIT_1B(256'hFFD9FFDD49FFD1357DE504C45DFFFFFFFD7FFFFD5FD5759C27FFFFFFFFFFDCD2),
    .INIT_1C(256'hFFD257D1D9FF3F9FFD85AC53FFFFFFFFFFFFFFFF5DD554C94CFFFFFFFFFFFF7D),
    .INIT_1D(256'hFFF17FD9FFFD1EFFFFF5EE755FFFFFFFFFFFFFFFFDF55D35709FFFFFFFFFFFF7),
    .INIT_1E(256'hDBF61FD1F7FED8DFFD7767657FFFFFFFFFFFFFFFF791592DB61FFFFFFFFFFFFF),
    .INIT_1F(256'h671EFD5BF7FDB79FFC56EBADFFFFFFFFFFFFFFFFD75450AB6647FFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n63,addra[14:13]}),
    .dia({open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,1'b0,open_n74}),
    .rsta(rsta),
    .doa({open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,inst_doa_i0_000}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF7D577CB81555555555617A055FA57DE977A8155555555555555555557DD5DD),
    .INIT_01(256'hFF77F50F97BFFFFFFFFF7F7A2DF4A97DE975A45FFFFFFFF557555555550D5FDD),
    .INIT_02(256'hFF477D7797DFFFFFFFFDB77A25DE995D615E115FFFFD75D588F556221F6AF793),
    .INIT_03(256'hFF475F6B347FFFFFFFFDE758B5F725FD617847F5FFF55C15C8DF415C1D5555DF),
    .INIT_04(256'hFF65F5D9B51FFFFFFFFDD758155A3A7D65D95FF5FFD7961DFD6D7C9557DDFEFF),
    .INIT_05(256'hFF65C7DA35DFFFFFD5F5D7505D7D21C5A569FFFFFFD7955565589F5FDFF59FFF),
    .INIT_06(256'hFF45F5D7577FFFFFD5F4DD6A5D6CAEB5A5AB7FFFFFDD55CB7889F5FFFDD73FFF),
    .INIT_07(256'hFF477DF727FFFFFFD5F515E275F02A5DADA97FFFFFF54DB80AFD7FFFFD547FFF),
    .INIT_08(256'hFF7779FD47FFD5FFD55DDFE155C32871A6A5FFFF7554528A8757FFFFFF65DE8F),
    .INIT_09(256'hFF5779FDA7FFFD7FD55F7DE3565A2A07AAAFFFFFD5BEAAA9D57FD7FFFF557723),
    .INIT_0A(256'hFF7547DD57FFFF5FD5DB7D417B1A6A80AA97FFF573A0AA7D7FF557FFFD75FFFD),
    .INIT_0B(256'hFFDD65DDDFFFD5D7D7DE7D7D59682AA82AB7F7F530A2A75FFFFD57FD7FD522FF),
    .INIT_0C(256'hFFDD7F5D5FFFF5AD7FDF7DBDE3BA320D6A57F5D7AAA9D55555557FFFFFDFBFFF),
    .INIT_0D(256'hFFD1565EB57F7B615F5575856D64B28D6AD7F57AAAA95555555F55FFFFF76FFF),
    .INIT_0E(256'h7FCF565EA557D4DA35575585AE8240AA6975D72AAAAAAAAAAAA297555FFDDBFF),
    .INIT_0F(256'h6FCD59F5AAD7D58CA5555777A5AB8CA9AB5F7EAAAAAAAAAAAAAAAA8757F758FF),
    .INIT_10(256'h4FF9D775AA9D55A02AC955759FA61C61AD576AA94AAAAAAAAAAAAAAA9D55D4FF),
    .INIT_11(256'h71755797AAA9D5EAAA31779EB8C176A1AD7AA58BF42AAAAAAAAAAAAAAA7575AB),
    .INIT_12(256'h17D45717AAAA9D52A955749E1E5CD54B85EC41D6E4AA554AAAAAAAAAAA09D559),
    .INIT_13(256'h35C7F475AAAAAA764BD5749418236E783D50D63F7F575F42A5CAAAAAA55575D7),
    .INIT_14(256'hED745D6D6AAAAAA0FFB5F67AC204142CF6F986D5A8DFD28AAFE9D555755555F7),
    .INIT_15(256'hF1D59DC5EAAAAA82243754DADA57B6245CD9AA10227FE76A808022F57FFD7FF5),
    .INIT_16(256'hF85595A96AAAA8285A175C411AA2AAA6120AAAAAAA8A3116AAAA80CA757FFFFF),
    .INIT_17(256'hFDDDD5895AAAAA9AFAB75E6BAAAAAAA80AAAAAAAAAAAA9326AAAAA8AA2D55FFF),
    .INIT_18(256'hFCF55DCA7AAAA9B51A4755EB6AAAAAAAAAAAAAAAAAAAA205E6AAAA80A20355F7),
    .INIT_19(256'hFF65F55A5AAAA9D929677D462AAAAAAAAAAAAAAAAAAAA9151CAAAAAAAA8B4D55),
    .INIT_1A(256'hFF57FD5A92AAAE02A947D5ACAAAAAAAAAAAAAAAAAAAAA89E62AAAAAAAAA81635),
    .INIT_1B(256'hFFF3FFDAB6AA892AA8D5D5A5AAAAAAAAAAAAAAAAAAAAAA4792AAAAAAAAAA8A59),
    .INIT_1C(256'hFFD757D686AA746AA8755732AAAAAAAAAAAAAAAAAAAAA94CF1AAAAAAAAAAAA0D),
    .INIT_1D(256'hBFFBFFD6AAAAD2EAAAF59592AAAAAAAAAAAAAAAAAAAAA86A244AAAAAAAAAAAA0),
    .INIT_1E(256'hD9FDDFDEAAA992CAAA579622AAAAAAAAAAAAAAAAAA26A79844CAAAAAAAAAAAAA),
    .INIT_1F(256'hDE1EDD5EAAAA5A4AA8751E0AAAAAAAAAAAAAAAAAAAA98968121AAAAAAAAAAAAA),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n122,addra[14:13]}),
    .dia({open_n126,open_n127,open_n128,open_n129,open_n130,open_n131,open_n132,1'b0,open_n133}),
    .rsta(rsta),
    .doa({open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,open_n154,open_n155,inst_doa_i0_001}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFC7FDBF77DFFFFFFFFFDFDFD7F761D77FDDFDFFFFFFFFFFFFFFFFFFFFFF557D),
    .INIT_01(256'hFFED5FFD765555555555E5DF575FB6D77FDDFBF55555555FFFFFFFFFFDD002F8),
    .INIT_02(256'hFFDDD7EF7EB555555557EDDF7F765C7777F76FF55557DFFDF5AAAB5D60B75FC7),
    .INIT_03(256'hFFDDF5F7DDB5555555579DDF5F78F4B777DD9D5F555FF76A97D57609D7FFFE1F),
    .INIT_04(256'hFFDF5F7F5DF5555555571DDDFFDBEF17775CB55F557D6BD7FF5AA9FFFD77F1FF),
    .INIT_05(256'hFFDF7D7DDF7555557F5D3DDD77C1559FF77C555555765FFF5827D5F5755F67FF),
    .INIT_06(256'hFFDF6F7E9DD555557F5FB7F5F76BFBCFF7FDD5555577FF7C0FDD5F55577E7FFF),
    .INIT_07(256'hFFDDC75F3D5555557F5EFF77DFAD754FF5FFD555555FFAE75FD7D55557D1FFFF),
    .INIT_08(256'hFFEDCF573D557F557FF47575FD36FD47F7F75555DFF7A7DFD5FD555555FA2B7D),
    .INIT_09(256'hFFEDE757DD5557D57FFCD755F59D7DD1FFF555557D69FFFD7FD57D5555FFD7D6),
    .INIT_0A(256'hFFCFDB77DD5555F57F76D75FDE5FBF79FFDD555FF675FF57D55FFD5557DF5555),
    .INIT_0B(256'hFFC7F37775557DFD7D79D76FDCBD5F797FDD5D5FEDF7F5F55557FD57D57457AA),
    .INIT_0C(256'hFFEFD9F5F5555FF7D57BD7E77C6FE7F27F7D5F7DFFFD7FFFFFFFD5555574FFFF),
    .INIT_0D(256'hFFEFF3F7DFD5DDFDF5F9DF5F7851EFF87F7D5FDFFFFD55555555FF55555DBFFF),
    .INIT_0E(256'hFFDBF9F7F7FD777F5FF9FFFFF3D555D67DDF7D7FFFFFFFFFFFFFD5FFF55767FF),
    .INIT_0F(256'hBFF3F6DDFF7D7DD5F7DBFDBDD9FEF9D4FDF5DFFFFFFFFFFFFFFFFFD5FD5DFDFF),
    .INIT_10(256'hDBDB74DDFFD7FFF57F77FD9DE975515CFFFD7FFD5FFFFFFFFFFFFFFFD7FF7D1F),
    .INIT_11(256'hFEF1FCFDFFFD7F7FFF6FDFF7E9AD08DEF7FFF5F60B7FFFFFFFFFFFFFFF5FDFE7),
    .INIT_12(256'h7FB9FE7DFFFFD7DFFD67DF77C083A2B6DFD17622B5FF555FFFFFFFFFFFFD7FDA),
    .INIT_13(256'h7F58DF9FFFFFFF57560FDFF54984B325DFA5096280A800B7F5DFFFFFF5555F7C),
    .INIT_14(256'hD7D2F5B77FFFFFF5824F5D5F354B8D41B6A8FF8AF500257FDA9D7FFFDFFFFF5F),
    .INIT_15(256'hD77CF7B77FFFFFDE9F4DFD5D35E3EDFA222755FFDD80957FFF555F5FD557D55F),
    .INIT_16(256'hF7FD7F5FFFFFFD7FA56DF5D6F555555F6DF5555555754857FFFFFD975FD55555),
    .INIT_17(256'hFE777FDDDFFFFFDD25EDF7FE55555557F555555555555C877FFFFFF55F7FF555),
    .INIT_18(256'hFFBFF75FDFFFFDE0759DFF76D55555555555555555555DDAB7FFFFD5FD5DFF5D),
    .INIT_19(256'hFFBF5FDF7FFFFE27D79DD75BD5555555555555555555540A0BFFFFFFFFF637FF),
    .INIT_1A(256'hFF4D57FFF7FFF09D57BD5FF35555555555555555555557CB7DFFFFFFFFFDCBDF),
    .INIT_1B(256'hFFE7557FD7FFD655571F5FDB5555555555555555555555F857FFFFFFFFFFDDA5),
    .INIT_1C(256'hFFF1FD77D7FF6BD5571F5D655555555555555555555557978DFFFFFFFFFFFF7A),
    .INIT_1D(256'hFFF6D577FFFF2F15551FDDED555555555555555555555715D15FFFFFFFFFFFF7),
    .INIT_1E(256'hA7FC7577FFFCA03555BDDFFD555555555555555555DD5CF7281FFFFFFFFFFFFF),
    .INIT_1F(256'hDA7DB7F7FFFF69F555BDD755555555555555555555677CFFC10FFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n181,addra[14:13]}),
    .dia({open_n185,open_n186,open_n187,open_n188,open_n189,open_n190,open_n191,1'b0,open_n192}),
    .rsta(rsta),
    .doa({open_n207,open_n208,open_n209,open_n210,open_n211,open_n212,open_n213,open_n214,inst_doa_i0_002}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFEBFFEC706FFFFFFFFF82F00FFF4BBFC3FF146FFFFFFFFFFFFFFFFFFFBEAFEE),
    .INIT_01(256'hFFEEAE1F6B3AAAAAAAABFBE41BE817AF92EB4DBEAAAAAAAFABAAAAAAAE1AEA3A),
    .INIT_02(256'hFF8AEBFE3AFBAAAAAAAB7AE55ABC73FFDEF8E2BBAAABEEEF15BAAA056AE0EB62),
    .INIT_03(256'hFF8AFAC768FAAAAAAAAA9BF16AAB5DAF9FF38AAFAAAFAC3E802F87BC7FABEEBF),
    .INIT_04(256'hFF9BAFBB3F6AAAAAAAAAFEE06AF070EEDBE5EAAFAABF6E7AFECAEC7EFFBBCDFF),
    .INIT_05(256'hFF9BCAB57EBAAAAABFAEFFF4FABA929A1B91FAAAAABB3FAEDEA56AFABAAE2FFF),
    .INIT_06(256'hFF8BBFBBAEEAAAAABFA9AFD0FB9C097F1E16EEAAAABBABCBA826AFAAABBF7FFF),
    .INIT_07(256'hFF9AEFA80EAAAAAABFAA6F90FEB1C5B21E46EAAAAABECFB4B06BFEAAABE9BFFF),
    .INIT_08(256'hFFFEA2AA9AAABFAABFFBFBD7FACE01F20C0FAAAAEFBCB5717FFFFEAAAACEBE12),
    .INIT_09(256'hFFFEA6AA5AAAAFEABFF3AF92F9F0100F011AAAAAAA3C5152AEFEAAAAAAFAE816),
    .INIT_0A(256'hFFBF8BBBEEAAABFBBFA7BF82E630C156057EAAAEC31E14EBFFFAAAAAABEEBEFE),
    .INIT_0B(256'hFFAFDAFBFFAAAF7EFFA8ABE3A7830455D42EAFFA23081EFEBAAAAAAAAABF52EA),
    .INIT_0C(256'hFFF3F3FBFAAABF4FAFA8EB7BC3302C4ED4BEAFFA1102FFFFFFFFEAAAAABB7FFF),
    .INIT_0D(256'hFFE2F8A86FEAF7D7FAEAEB5FD987205B90FEAAA40012EAAAABEEFFFBAAAEDFFF),
    .INIT_0E(256'hFFCEE9A94AFFBDF1FFFAEF9A4930D30582AFBFC45401414001546FBFFAABA3FF),
    .INIT_0F(256'h9FCEE3EB55FEBE7A1AAAFE9E0F021F0242FAE045501500000005543ABFAAF9FF),
    .INIT_10(256'hDEF3FBEF002BEA4A8186BEAE6A4C388703EB8517A4010105400000552EFFB8EF),
    .INIT_11(256'hB6BAFF3E0003FFC540F3ACA834C3BD064BE41B06B88000000000005051FFFE17),
    .INIT_12(256'h28F8BB3F01052AE553FBFC6829F8BF873B9ED7B89B05BEE0555001554556BFA6),
    .INIT_13(256'h4ACAB8BE415541BDE6ABE97B7016EBE02BA9B95ABEBFAE884F3000005EBFAFBF),
    .INIT_14(256'hDFE9FFCBD015404FFE7EE8A09058304DBD32D67EF4BEF4500EC2EAAAABFFFFEE),
    .INIT_15(256'hE7BF6FDFD0014025546AADA4C57D912DEDA0150000BBDE94111054EFFFFEEABF),
    .INIT_16(256'hF1AB2A56800002D1B02BA9FAC5515112344555555505663D000045C1EFEEAAAA),
    .INIT_17(256'hFBFBBB13E4001574D0ABA8C1555414515555555555555A358400005401BFAAAA),
    .INIT_18(256'hFDEFEB80A400133A148BBB8415555551555555555555541A9C00042A0016EEAE),
    .INIT_19(256'hFF9BAFE5E40003E1548ABABE15555555555555555541526EA800000000065AFF),
    .INIT_1A(256'hFFBFAFE03D00195555CFAE4C5555555555555555555551A9C540000010031F2F),
    .INIT_1B(256'hFFE6BEE57900271555EFFF1855555555555555555555500E38000000140030F6),
    .INIT_1C(256'hFFEBFEBD6900E95555FFFFA45555555555555555555555D0E6000000000000CE),
    .INIT_1D(256'h3FF3EAB95401A7D554EF7E655555555555555555555555C048A000000000000D),
    .INIT_1E(256'hA7FBFAB95006248555BE6D31555555555555555555C153C1D8F0000000000000),
    .INIT_1F(256'hB93DBBFD5005B00555AF6D01555555555555555555401A2C79E4000000000004),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n240,addra[14:13]}),
    .dia({open_n244,open_n245,open_n246,open_n247,open_n248,open_n249,open_n250,1'b0,open_n251}),
    .rsta(rsta),
    .doa({open_n266,open_n267,open_n268,open_n269,open_n270,open_n271,open_n272,open_n273,inst_doa_i0_003}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF9AAB3FFABAAAAAAAAAFBBFAAABD2EAFEABEEBAAAAAAAAAAAAAAAAAAAFFBAFF),
    .INIT_01(256'hFF9AABAFFDFAAAAAAAAA9ABBBEAF78EAEEABB2EAAAAAAAAAFFFFFFFFFBE110A1),
    .INIT_02(256'hFFAEAA9BAD6AAAAAAAAADEBAFAADFCAAAEAFCBAAAAAAABFBAE1554EB900AEFCB),
    .INIT_03(256'hFFBEAABFAF3AAAAAAAAB3EAFBAB1AF7AAEBF3EAAAAAAFFD13BBFF857AEFEB96F),
    .INIT_04(256'hFFBEAAA2BABAAAAAAAAB6AAEAAA78F3AEAAF3AAAAAABD0ABFFA117EFAAAAE7FF),
    .INIT_05(256'hFFBEEEAFBAAAAAAAAAAB6ABAAAD6EA6EEAEFEAAAAAADABFFB00BAEAAAAABCFFF),
    .INIT_06(256'hFFBE9AAD7AAAAAAAAAAE3ABFAA92F69BEAEBAAAAAAAAFEF142FEEAAAAAA9BFFF),
    .INIT_07(256'hFFAE8EAE6AAAAAAAAAADBABBAA4BFE8AEABEAAAAAAABB41AFFFAAAAAAAB2FFFF),
    .INIT_08(256'hFF9ACBAB6EAAAAAAAAA8EAEEAA2DBFDAFFFAAAAAAAEA4AFEBBAAAAAAAAA104EB),
    .INIT_09(256'hFF8ADFABFEAAAAAAAAA9EAFAAF7FBFA3FEFAAAAABF97BEAEEAAAAAAAAAAFAEF8),
    .INIT_0A(256'hFFDAF7AABAAAABAAAABDEAEAADBF3EA2FAAAAAAAA9EFEBFAAAAAAAAAAAABBFFF),
    .INIT_0B(256'hFFDEB7AAAAAAAAEAAAB2EA9AAC3FBFA2EBEAAAAB9BFFFAAAAAAAAAAAAAA8BC55),
    .INIT_0C(256'hFFCAB3AAAAAABAFEAAB6AADAF9CF9FE0EBAAAAABFEFEEAAAAAAAAAAAAAA9FFFF),
    .INIT_0D(256'hFFCBA6EBEAAABFBAAAB7AAEAB7BFDBB4AFEAAABFFFEEAAAAAABEAAAAAAAA3FFF),
    .INIT_0E(256'hBFE7B7EBBAAAAABEFAA6AA2EF6FBEBF9BEAAABFBABFEBEBFFEABEBAAAAAA9BFF),
    .INIT_0F(256'h7FE7B8EBABEAAABBEAF7AA6BF7FDE3FCFFAAABBAAFEAFFFFFFFAABFBAAAAA2FF),
    .INIT_10(256'hA7F2ADAAFFEAAAFFFFBFAB6AC3EEB6BCFAAEFAFFBAFEFEFABFFFFFAAEEAAAF7F),
    .INIT_11(256'hF9B2A9ABFFFEEAFABFDEAA3BC24A11FDBEBFEFE943FFFFFFFFFFFFAFAFBAABDF),
    .INIT_12(256'hFE67EDABFEFAEEBAAFDEABFF85425028BAE3E8016BFFBEFFAAAFFEAABAAFAAF4),
    .INIT_13(256'hAFF4EF7AFEAABFBEFD4AAEEB8209055EBE0F57C05441013FBFFFFFFFFEAAEAA9),
    .INIT_14(256'hFEA4AB2AAFEABFBF158AAEEF2F824AC7791038414F504EBFF17EEAAAAAAAAAAB),
    .INIT_15(256'hFAA8FA6AEFFEBFF92ADEABBB2F821B84110ABFAAAB547EABEBEABAEAAAAAAAAA),
    .INIT_16(256'hFEEEBBFEBFFFFFAF1EDEABBC6FFBEFF8DFEFFFFFFFAE90BEFFFFAE6BAAAAAAAA),
    .INIT_17(256'hFCEAAAAEABFFEABF5E0EAABCBFFFFFFFFFFFFFFFFFFFE05BBBFFFFBFFBEAAAAA),
    .INIT_18(256'hFE7AAAAFBBFFEFD4BE7EAAF9BFFFFFFFFFFFFFFFFFFFFEB46FFFFBFFFBABBAAA),
    .INIT_19(256'hFF3EAAAAABFFF84BFE2EBAB0BFFFFFFFFFFFFFFFFFFFFC5046FFFFFFFFE9EFAA),
    .INIT_1A(256'hFFCAAAAFFEFFE56BFF7ABAF7FFFFFFFFFFFFFFFFFFFFFF06FEBFFFFFEFFFB1EA),
    .INIT_1B(256'hFFDBAAAEAAFFEDFFFF7AEBF2FFFFFFFFFFFFFFFFFFFFFFB0BFFFFFFFEBFFFF0F),
    .INIT_1C(256'hFFE3AAAEBAFFC3BFFF3AAACEFFFFFFFFFFFFFFFFFFFFFF7B0AFFFFFFFFFFFFE4),
    .INIT_1D(256'hBFFDEAAAAFFE583FFF2AEA8FFFFFFFFFFFFFFFFFFFFFFE3FE6BFFFFFFFFFFFFE),
    .INIT_1E(256'h0EFCEAAEAFF8443FFE6AAB9BFFFFFFFFFFFFFFFFFF6BF92F103FFFFFFFFFFFFF),
    .INIT_1F(256'hE5AF3AAEAFFA82BFFF7BAFFBFFFFFFFFFFFFFFFFFFDAF092934BFFFFFFFFFFFB),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n299,addra[14:13]}),
    .dia({open_n303,open_n304,open_n305,open_n306,open_n307,open_n308,open_n309,1'b0,open_n310}),
    .rsta(rsta),
    .doa({open_n325,open_n326,open_n327,open_n328,open_n329,open_n330,open_n331,open_n332,inst_doa_i0_004}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFE5F67FB5E77FFFFFFF4D4D435532FD37545C7FFFFFFFFFDFF575FFFD7F4234),
    .INIT_01(256'hFFF5FDDE932F7FFFFFF777C501D7D3D5957DDD75FFFFFD5DF75FFD755CEE2638),
    .INIT_02(256'hFFEDDFD75FDF7FFFFFF575457FD1941D9FD1FDF5FFDFF7FCBABF54969546B76B),
    .INIT_03(256'hFFE5F7F3F4FFFFFFFFF5A76E07DED7FDBFEFCF55FFFD59172F02938C43FDFDAF),
    .INIT_04(256'hFFE7FF7146DFFFFFFFFF854CFFC7F7275BC57FF5FFF4BCEDFF1B54F77D77C277),
    .INIT_05(256'hFFE73DFE6F7FFFFFFFF6BF5CBF6ACACF511F97FFFFD1E5DD0EB8417F7D5D93FF),
    .INIT_06(256'hFFC7F7F7C7FFFFFFFFFDBFF275355F4C5B7EFFFFFFF7579291FEB7FFFF759FFF),
    .INIT_07(256'hFFC551FCAFFFFFFFFFF57FF9FFF5DA8370F57FFFFFD75519F547FFFFFF685FFF),
    .INIT_08(256'hFF555BFD35FFFF7FFFF4B7367C3D756B5759FFFFFD5B73F77A7DFFFFFFE7F492),
    .INIT_09(256'hFFD7F9F745FFDDFFFFD05FA352163460FFFFFFFFF47C775E37D57FFFFFFF70CA),
    .INIT_0A(256'hFFCF4F774FFFF47FFFF37D2D5F1DFD16FF45FFFD4B9DD765DFD7FFFFFFF54AA8),
    .INIT_0B(256'hFFC97B7FD7FFF455D55B5F13E4DF8D1EFFD5F5F7F77D53DFFDF7DFFFFFDA2075),
    .INIT_0C(256'hFFF3C0F655FFC5F9D5DE7DFDB4BD5D117D9FFFDE5FFE1D555557D7FFFFF67FFF),
    .INIT_0D(256'hD7FDD8F757FFEE5657F45D0D9FAF75EEB73FD7EFFFF682AA8801D7F7FFF57FFF),
    .INIT_0E(256'h77C7D675717F5387C5F5DF17537A63EB3CFFF4DFFFD555555555E2F5FFFD57F7),
    .INIT_0F(256'hDFF9F5F5F7BDFCFBDBE5FF6EC957D760F67F5B7FFFFFDFFFFFFF55F2D7FD50FF),
    .INIT_10(256'h4DEBD2547D6FFDDF55D9FE54F61F98A8F3D7BFDD37FFFFFFFFFDD755E3FFF40D),
    .INIT_11(256'hD570F496F5D4959DFFD7D61D5CD40C40F3F57553A6FFFFFFFFFFFFFFD725FD73),
    .INIT_12(256'h9CDEF516F57DCBE55DC15531CAADF973FD63D3F97BF73E5FFFFFFFFFF5D6FF45),
    .INIT_13(256'h8F27FFE777FFD5AF510F7F5B835454B045DF898449FCA2C7F577D75FF6821FD4),
    .INIT_14(256'h69737EE71FFFFF5FC65FFFB56468F6F9F33BCD1037C7342F4FC69DFFFDF57FDD),
    .INIT_15(256'hCB5C7F5B1FFFFF7DDF77FCE6724766F5BFE1EADFD6BF44BFF6802EB55F7FDFFF),
    .INIT_16(256'hF35CD50F7FFFF7F6F9F5F47F1AA22A8562B2AAAAAAF0DE3575557A65B5FFFFFF),
    .INIT_17(256'hF59FF586E7FFFFDE8165F6F4AA828AAAAAAAAAAAAAAA2D619FFFF5C2279DFFFF),
    .INIT_18(256'hFF7FD76767FFF5F3CBA5FFBA6AAAAAAAAAAAAAAAAAAAA8ADF5FFFFFDD4AED77F),
    .INIT_19(256'hFF57FFC537FFDD20A935E7BDEAAAAAAAAAAAAAAAAAAAABA7457FFFFFD55BD17F),
    .INIT_1A(256'hF7AFFFDF47FFFA7CA8DFE75AAAAAAAAAAAAAAAAAAAAAA0777ADFFFFFFFF57DF5),
    .INIT_1B(256'hFFD9FFF749FFE948AA478661AAAAAAAAAAAAAAAAAAAAA8C99DDFFFFFFFFFF6F2),
    .INIT_1C(256'hDFF87FF7F1FD6ACAA8CF046FAAAAAAAAAAAAAAAAAAAAA83E947FFFFFFFFFFD75),
    .INIT_1D(256'hBFF9DFF1FFF71BAAAA5FCEC0AAAAAAAAAAAAAAAAAAAAA0E080BFFFFFFFFFFFFF),
    .INIT_1E(256'h9BF69FF1FFDEDB0AAADD4F4EAAAAAAAAAAAAAAAAA804A5D874B7FFFFFFFFFFFF),
    .INIT_1F(256'hE51EB7FBFFFD986AABD649B6AAAAAAAAAAAAAAAAA2612DFF28CDFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n358,addra[14:13]}),
    .dia({open_n362,open_n363,open_n364,open_n365,open_n366,open_n367,open_n368,1'b0,open_n369}),
    .rsta(rsta),
    .doa({open_n384,open_n385,open_n386,open_n387,open_n388,open_n389,open_n390,open_n391,inst_doa_i0_005}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFD75FDEB03DD555555541D28FFF87D749FDA8B555555555755FDF5557575DFD),
    .INIT_01(256'hFF5D552F151555555555F572AF542B5749542E5555555557F55FFD755587F679),
    .INIT_02(256'hFF4D557D3D7555555557B5D0657C8BF7C974915555555F75C09FF48815C35791),
    .INIT_03(256'hFF6555CB945555555555A5F21D778357697245555557549FAA5DC9D49DFF757F),
    .INIT_04(256'hFF4575733D15555555577DF295F098DD055BD555555FB41F7FCBDE17D5555CFF),
    .INIT_05(256'hFF45CD7895555555555F75C8D57581658F43F5555577BDD7E55815D555551FFF),
    .INIT_06(256'hFF45DD55DD555555555E95685766A6BD8D89D55555555543D0295D55557FBFFF),
    .INIT_07(256'hFF65DF5DBD5555555555B5E05579AA752709D555555FCF3AAA15555555F67FFF),
    .INIT_08(256'hFFFD5F5545555555555755E7D54B8931008F5555577C5AA82FD5555555FD7C25),
    .INIT_09(256'hFFFD5157A555575555775569F6482A0F800D5555753C2801DD5555555577F5A2),
    .INIT_0A(256'hFFF54D55D55557D555795743D980C02B003D5555D30A001755555555555D7555),
    .INIT_0B(256'hFF57CF5575555F3D555855D55B622A0A801D55571A802F7555555555557F80D5),
    .INIT_0C(256'hFFD77757F5557F8F5555D71FC332BA27007555752001FFFFFFFD55555557BFFF),
    .INIT_0D(256'hFFD17FD49D555BE3F575D7AFE74E9AA748D55558000BFD5557DD7D55555DEFFF),
    .INIT_0E(256'hFFCD54560DD57EDABF555525AEA02A0A41555F80002800000000975F555753FF),
    .INIT_0F(256'hEFC5735C005555A405F5575D2CA9268981D5D400000000000000002D7D55F2FF),
    .INIT_10(256'hC5DD75DF001D550002C1575F9F82264B055DC02862000000000228001D5554DF),
    .INIT_11(256'hD375DFFD0A03FFC200B35D1698EB7CAB05580001FE0000000000000002FF550B),
    .INIT_12(256'h9D7E573F0A8015D2A8175C94345E7741A76621F4660A412000000000008BD559),
    .INIT_13(256'h9FEF5CDD8800027029555C963C0BEEDA9759DA9EF7575D68202800AAA17D557F),
    .INIT_14(256'hEFF4D577C000000ADE9D5CDAF981158D7C5FB6D22257F6008DE1D555575FD555),
    .INIT_15(256'hDB77B76FC0000002871554D8DD4FB5E4764DD5DFFF95E3402220AB5FF5555555),
    .INIT_16(256'hFA5F95A9E000000A773554E91555F576ADFD555555FD11828AAA0AC2FF555555),
    .INIT_17(256'hF7F5D7EBD000000877A55741D57D7557F55555555555F19A60000A88007F5555),
    .INIT_18(256'hFED555C8D000083D17A55749555555555555555555555DED620000020029DD55),
    .INIT_19(256'hFF655550500029CDD5255566D5555555555555555555579D9E8000000AA9EDD5),
    .INIT_1A(256'hFFFD55509800262D55CDFD85555555555555555555555F960A200000000A3D3F),
    .INIT_1B(256'hFFD95558140033B557DD7F8155555555555555555555577B0A000000000028D9),
    .INIT_1C(256'hFFD7D5502C02235557F5FDAB5555555555555555555555A7390000000000028F),
    .INIT_1D(256'hFFF3555C080A76955555BD2D555555555555555555F55FDFFC4000000000000A),
    .INIT_1E(256'h9BF77554002118B55775362D55555555555555555735559FC6E8000000000000),
    .INIT_1F(256'h763E955C00007555565D3EAD5555555555555555553D71C3DE92000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n417,addra[14:13]}),
    .dia({open_n421,open_n422,open_n423,open_n424,open_n425,open_n426,open_n427,1'b0,open_n428}),
    .rsta(rsta),
    .doa({open_n443,open_n444,open_n445,open_n446,open_n447,open_n448,open_n449,open_n450,inst_doa_i0_006}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFF65573DF55555555555F75F5557E1557D55FD55555555555555555555FD75DF),
    .INIT_01(256'hFF65575FFEF555555555657F7D5FB4D5FD55F1D5555555555FF557DFF750035E),
    .INIT_02(256'hFF555567569555555555ED7F355EDC557D5FC755555555D7DDE009576017DFC7),
    .INIT_03(256'hFF5D557F5F3555555557FD5FF57276B55D7F3D555555FF60DD7F742B5D55569F),
    .INIT_04(256'hFF7D7555757555555555955D555B6F35755E35555557C15DFD5C29DD5555DBFF),
    .INIT_05(256'hFF7DD55F755555555555955555E9F59DF5FED555555ED77D7005DD555557CFFF),
    .INIT_06(256'hFF7DE55E355555555555F57F5569F965F5F755555555FDF605FDD55555567FFF),
    .INIT_07(256'hFF5D4D5535555555555E55F75584FD45DDFD555555557865FF7555555551FFFF),
    .INIT_08(256'hFF65CD579D5555555554D5D1559E7C65F7F5555555D585FFF7555555557209D7),
    .INIT_09(256'hFF45EF55FD5555555556D5F55F1F7F537FFD55555F6BFFFDD5555555555D7D77),
    .INIT_0A(256'hFF65F35575555755555ED5D55E5F3FD3FFD5555556FFFF755555555555577FFF),
    .INIT_0B(256'hFFED715555555555557DD5655C3F7FF1FFD5555567FFF7555555555555547DAA),
    .INIT_0C(256'hFFC57355555575FD557955EDF6CF6F587F555557FFFDD555555555555556FFFF),
    .INIT_0D(256'hFFC75357D5557F7D555B55D57A7BE7787FD5557FFFFD5555557D555555553FFF),
    .INIT_0E(256'h7FDB7BD7F555555DF559555DF9F757F67D5557FFFFFFFFFFFFFFDF55555567FF),
    .INIT_0F(256'h3FDB54D5FFD55577F55B5797F9FEDBFCFF5557FFFFFFFFFFFFFFFFF7555555FF),
    .INIT_10(256'h5BF95E55FFDD55FFFFFF5595C1F7597CF5557FFD7DFFFFFFFFFFFFFFDD555FBF),
    .INIT_11(256'h747156D7FFFDD5FFFFED5577E18520FEFD7FF5DE03FFFFFFFFFFFFFFFF7557EF),
    .INIT_12(256'h7591DE57FFFFDD7FFD4D57FF4A09801E75DB548297FF557FFFFFFFFFFF7DD5F8),
    .INIT_13(256'h55D2D735FFFFFF777E8555F74B0E192D7D0C2D4B2A02023FF57FFFFFF555D556),
    .INIT_14(256'hFD7857357FFFFFFF23C5575FBFCF25E8B628752F572281DFF2BDD55555555557),
    .INIT_15(256'hF554D595FFFFFFF6174D57FF9F7947D800B5FFDFFDC0B57FD7D577D555555555),
    .INIT_16(256'hFDD5F7FD7FFFFFFF0FCD577C5FF7DFF5FFFFFFFFFFFFC057FFFFDD9775555555),
    .INIT_17(256'hFCD5D5DD5FFFFFDF8F7D577C7FFFFFFFFFFFFFFFFFFFD6277FFFFF5FF7D55555),
    .INIT_18(256'hFDB555DF7FFFFDE2DFDD55F47FFFFFFFFFFFFFFFFFFFFF5097FFFFFFF7577555),
    .INIT_19(256'hFF3D555FDFFFF6B5FDFD7571FFFFFFFFFFFFFFFFFFFFFC0089FFFFFFFFD69F55),
    .INIT_1A(256'hFF45555FDFFFDA9FFD35D5FBFFFFFFFFFFFFFFFFFFFFFF697DFFFFFFFFFF60F5),
    .INIT_1B(256'hFFE7555FF7FFFCFFFF35D7FDFFFFFFFFFFFFFFFFFFFFFF7E5FFFFFFFFFFFFF0F),
    .INIT_1C(256'hFFD35557F7FF7F7FFFB557FFFFFFFFFFFFFFFFFFFFFFFDF7E5FFFFFFFFFFFFD8),
    .INIT_1D(256'hFFFED557FFFD8D7FFF15D5FFFFFFFFFFFFFFFFFFFFFFFD3FD17FFFFFFFFFFFFD),
    .INIT_1E(256'hCDFCD55FFFFC827FFD15D75FFFFFFFFFFFFFFFFFFF57F457A03FFFFFFFFFFFFF),
    .INIT_1F(256'hDA5FF55FFFFF4B7FFF37DF7FFFFFFFFFFFFFFFFFFF65F677EB8FFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_000000_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n476,addra[14:13]}),
    .dia({open_n480,open_n481,open_n482,open_n483,open_n484,open_n485,open_n486,1'b0,open_n487}),
    .rsta(rsta),
    .doa({open_n502,open_n503,open_n504,open_n505,open_n506,open_n507,open_n508,open_n509,inst_doa_i0_007}));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hDE7F7657FFFD5F5FFE54E977FFFFFFFFFFFFFFFFD5E51567CE23FFFFFFFFFFFF),
    .INIT_01(256'h7DE574967FFCC97D76F44B5FFFFFFFFFFFFFFFFFDD1708675927FFFFFFFFFFFF),
    .INIT_02(256'hFF5C16147FFF6D7D77B7769FFFFFFFFFFFFFFFFFDFB3E26D7E8FFFFFFFFFFFCF),
    .INIT_03(256'hFF5DC5EC7FF5ED7D73D9F53FFFFFFFFFFFFFFFFFD7F3BD5D7765F5FFFFFFFD1A),
    .INIT_04(256'h0555DD9E7FCA6FFD70D184DFFFFFFFFFFFFFFFFFD5F3B8B5D528B5FFFFFFFFEA),
    .INIT_05(256'hD9597D99FFFD3FDD767BCF5FFFFFFFFFFFFFFFFFD5F2F5D7D5566FFFFFFFFF45),
    .INIT_06(256'hE75D5F751F947FFF5493F81FFFFFFFFFFFFFFFFFD5F3A9FDD5D8F3FFFFFFFF74),
    .INIT_07(256'hF4D97F6C9D59D7F7DC9F9CBFFFFFFFFFFFFFFFFFFFDEC9F75750F9FFFF7C3FFF),
    .INIT_08(256'hFF7E27453FD97D5FDC5DB847FFFFFFFFFFFFFFFFFFDFD77753F677FFFFF9D3FF),
    .INIT_09(256'hFD6709DD7D197FFFFCE7F60DFFFFFFFFFFFFFFFFFFDFAF74308D7DFFFFFD95BF),
    .INIT_0A(256'hFF6D8C59FDBFFFD5F14CC52FFFFFFFFFFFFFFFFFFFDF5FAE5FD1CEFFFFFD36F9),
    .INIT_0B(256'hFDD76C317D07FCD859EF8A185FFFFFFFFFFFFFFFFFDFF633757DB1BFFFF5C3E8),
    .INIT_0C(256'hFFFDF7AFF10F7778F8E6ADE557FFFFFFFFFFFFFFFFFFD965DFFFDE9FFFFFF2F7),
    .INIT_0D(256'hFFF877DAF78F7055D6E43B0F957FFFFFFFFFFFFFFFF5EDDFFFFFD0DFFFFFD6BD),
    .INIT_0E(256'hFFF69D3EF7BDEC250B00F157A77FFFFFFFFFFFFFFFF54345FFD7CAFFFFFFDD2F),
    .INIT_0F(256'hFFFF51DFFE5F8002408ECF9DDF7FFFFFFFFFFFFFFDDF2795FFD7746FFFFFFDFF),
    .INIT_10(256'hFFFFEDBABE5FA296C2C5C8D1737FFFFFFFFFFFFFFD7433557FD758B77FFFFF6B),
    .INIT_11(256'hFFFF8D4E6657003DF9EE7388D0FFDFFFFFFFFFFFD53AF77FFFD7DF57FFFFFFC8),
    .INIT_12(256'hFFFFE2D1847501D541770498E5DFF77FFFFFFFFFD42977FFFFFFD7C7FFFFFFF9),
    .INIT_13(256'hFFFFDCE8DB37235FF1E821AA9995F77FFFFFFFFD5A2DFFD57FFFDF29FFFFFFFC),
    .INIT_14(256'hFFFFF8B70D97AFFFF3875C18AD15FF57F5FFFFFD679DDFF5F5F7FE1FFFFFFFFF),
    .INIT_15(256'hFFFFFE7C009F9BFFF91E50426DBD7DFFFFFFFFF79CC3D555FDD7FF37FFFFFFFF),
    .INIT_16(256'hFFFFFD137E5F97FFF719FF34F5B17557FDFFFFDD69EFF0727757FF73FFFFFFFF),
    .INIT_17(256'hFFFFFF9FA8751FFFF4CEFFF1AAD57A5D757FDF758C5ADFFD50AF5FE55D5FFFFF),
    .INIT_18(256'hFFFFFFF6053703FFFEA7FF6F14CA74DDDF7FD57ADA3E28160BD75F24EFFFFFFF),
    .INIT_19(256'hFFFFFFE8DF8F2BFFFF5FFCC3D53B3DDD657FF5CC4EE0000B36BD7F1A435FFFFF),
    .INIT_1A(256'hFFFFFFF892EF0BFFFC8FFC3EFD8EF95F735FF6394000962E03E77F50CB2FFFFF),
    .INIT_1B(256'hFFFFFFE255ED23FFFD5FFFFDFC06365FCFDD71300C4DFFFF1C31D57E8BFFFFFF),
    .INIT_1C(256'hFFFFFFC321355FFFFDFFFBF77F85E0FFEF570B4C30235555DE82D571461FFFFF),
    .INIT_1D(256'hFFFFFFE20CF55FFFFFAFFA1EFF37E1FF995FDB222FFFF55EB785DF915F47FFFF),
    .INIT_1E(256'hFFFFFFE1A51D63FFFF5FF29A7F56995791DF7A179BFFFFFFD52BFFF7EFC7FFFF),
    .INIT_1F(256'hFFFFFFDD8BFDDFFFFF9FF1227FEBF155D38534F35BFFFFFFFA27F5458707FFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n535,addra[14:13]}),
    .dia({open_n539,open_n540,open_n541,open_n542,open_n543,open_n544,open_n545,1'b0,open_n546}),
    .rsta(rsta),
    .doa({open_n561,open_n562,open_n563,open_n564,open_n565,open_n566,open_n567,open_n568,inst_doa_i1_000}));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hD54F7756AAA8C2AAAA7516EAAAAAAAAAAAAAAAAAA8E2E0121FCAAAAAAAAAAAAA),
    .INIT_01(256'h7D568FD7AAA966AAA2D5944AAAAAAAAAAAAAAAAAA8381B62A5D2AAAAAAAAAAAA),
    .INIT_02(256'h7F55DF55AAA85AAAA116A00AAAAAAAAAAAAAAAAAAA70ECDAA9BAAAAAAAAAAA9A),
    .INIT_03(256'h1F5D75B7AAA19AAAA7BEA12AAAAAAAAAAAAAAAAAAA866B8AAA14AAAAAAAAA810),
    .INIT_04(256'h1555DD67AA92AAAAA73E83AAAAAAAAAAAAAAAAAAAA83626AAA536AAAAAAAAA98),
    .INIT_05(256'h7D557DE5AAA56AAAA196E32AAAAAAAAAAAAAAAAAAAA5ACAAAA01DAAAAAAAAA1D),
    .INIT_06(256'hDD5A5F696A732AAAA156426AAAAAAAAAAAAAAAAAAAA580AAAA89F6AAAAAAAA22),
    .INIT_07(256'hF0559F51689CAAAAA9DAC56AAAAAAAAAAAAAAAAAAAA840AA02A6F8AAAAA96AAA),
    .INIT_08(256'hFD97F77A6AB0AAAAA95AE45AAAAAAAAAAAAAAAAAAAA8E282A8A97AAAAAAAE6AA),
    .INIT_09(256'hFD75B5DAA896AAAAA378410AAAAAAAAAAAAAAAAAAAA85AAB322060AAAAAADE6A),
    .INIT_0A(256'hFFA54756A8CAAA80A1FAC5EAAAAAAAAAAAAAAAAAAAA8CA4C4A8A29AAAAAA4344),
    .INIT_0B(256'hFFF944DE289AA87083DB19F9AAAAAAAAAAAAAAAAAAAAA9192AAA736AAAA01F3C),
    .INIT_0C(256'hFFFD47B6A75AAA8AD6D39ABE2AAAAAAAAAAAAAAAAAAAA74CAAAA898AAAAA85F2),
    .INIT_0D(256'hFFF2FFCDA25AA500AC99B4656AAAAAAAAAAAAAAAAAAA97D2AAAA870AAAAA817F),
    .INIT_0E(256'hFFFFD9B9A1AA8E087B39DE8798AAAAAAAAAAAAAAAAAA335AAAAA94AAAAAAA8FF),
    .INIT_0F(256'hFFFCF46AABAA50003CB75C4348AAAAAAAAAAAAAAAAAA6D6AAAAAA8DAAAAAA817),
    .INIT_10(256'hFFFFFEB5612A51350015794FDEAAAAAAAAAAAAAAAAA912AAAAAAA5A2AAAAAA2D),
    .INIT_11(256'hFFFF7607D12A52688F194E1B71AAAAAAAAAAAAAAAA4CE0AAAAAAA822AAAAAA93),
    .INIT_12(256'hFFFFC986DB0A50AA9BA92D6744AAAAAAAAAAAAAAA91B2AAAAAAAAA02AAAAAAA5),
    .INIT_13(256'hFFFFF58B834A79FFF7AFE096CB6AAAAAAAAAAAAAA6E482AAAAAAAAB6AAAAAAA9),
    .INIT_14(256'hFFFFF45C696A73FFFE4E8823570AA8AAAAAAAAAA9FBA2AAAAAAAA9CAAAAAAAAA),
    .INIT_15(256'hFFFFFE17556A67FFFEFFD4013CCAABAAAAAAAAAA56F68000AAAAAA3AAAAAAAAA),
    .INIT_16(256'hFFFFFF10232A67FFF653FD70AB9EA32AAAAAAAA842700DF20A0AAA96AAAAAAAA),
    .INIT_17(256'hFFFFFF60B7AA6FFFFF32FFFF8818A82AAAAAAAA383F22AA0022AAA92880AAAAA),
    .INIT_18(256'hFFFFFFD1512A73FFFE35FF5F7155A4AAAEAAAA26DFC82821F61AAA585A2AAAAA),
    .INIT_19(256'hFFFFFFE8211A73FFFEDFFFEBDAA166AA04AAA810EF800002596AAA7A5C8AAAAA),
    .INIT_1A(256'hFFFFFFF85E5A53FFFFCFFC31F715A4AA12AAA0EE0001D7D00052AA1279DAAAAA),
    .INIT_1B(256'hFFFFFFEAE2DA53FFFD8FF73CFF83EDAA9AAAA36009E2AAA89000AA1C86AAAAAA),
    .INIT_1C(256'hFFFFFFCB96CA3FFFFF2FFF3EFF6359AA12AAE20307D6AAAA8A85AA1B594AAAAA),
    .INIT_1D(256'hFFFFFFC2224A1FFFFF7FF6BE7F0960AAB6A8CAE77FFFFFF74808AAD3A9E2AAAA),
    .INIT_1E(256'hFFFFFFC386CA27FFFF5FF62EFF4E58AA1689165537FFFFFFD936AA919D62AAAA),
    .INIT_1F(256'hFFFFFFF383AAA1FFFF7FF782FFDDD0A8564E53F1D3FFFFFFFD22AA2140A2AAAA),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n594,addra[14:13]}),
    .dia({open_n598,open_n599,open_n600,open_n601,open_n602,open_n603,open_n604,1'b0,open_n605}),
    .rsta(rsta),
    .doa({open_n620,open_n621,open_n622,open_n623,open_n624,open_n625,open_n626,open_n627,inst_doa_i1_001}));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7DA99DFFFFFDAD5557BDD79555555555555555555739DBCD7057FFFFFFFFFFFF),
    .INIT_01(256'hD7DABD7FFFFDBD555FBDD7B5555555555555555557464FBD5E17FFFFFFFFFFFF),
    .INIT_02(256'hD5FD2D7DFFFFB5555E7FF5F5555555555555555555C73D3557CFFFFFFFFFFFDF),
    .INIT_03(256'hF5F7DFDDFFF675555C77F65555555555555555555571D47555C9FFFFFFFFFD65),
    .INIT_04(256'h5FFF777DFFD775555CF7745555555555555555555574DFD555C07FFFFFFFFFC1),
    .INIT_05(256'hE7F7D777FFFA15555CF79CD55555555555555555555C535555F89FFFFFFFFF5A),
    .INIT_06(256'hDBF7F5FF7F6AD5555C77B7D55555555555555555555EDF55557CA7FFFFFFFF75),
    .INIT_07(256'hFDF6F5DD7DEB5555547F18D5555555555555555555559F55FD5F25FFFFFD7FFF),
    .INIT_08(256'hFEFF3DDF7FE7555554FF31B555555555555555555555155D5D57AFFFFFF6B7FF),
    .INIT_09(256'hFF9F477FFD6D555554DFB85555555555555555555555355447F7ADFFFFFEAB7F),
    .INIT_0A(256'hFFFF59F7FD15557F56DD9A355555555555555555555535D1B55D49FFFFFF3CB5),
    .INIT_0B(256'hFFEFD9777FF5550D76DE6F2F555555555555555555555766D555C27FFFF5C7C3),
    .INIT_0C(256'hFFD3FA5FF635555F01D44549D55555555555555555555E9B5555785FFFFFF1FE),
    .INIT_0D(256'hFFF5DAB5F6355FFF51DC4DFAD55555555555555555557AAD555570DFFFFFDC7F),
    .INIT_0E(256'hFFFC7E6DF6D57357FE54AD7AF5555555555555555555C6B5555570FFFFFFFF1F),
    .INIT_0F(256'hFFFFB7BFFC55C000815881F6B55555555555555555553AD55555549FFFFFFDEF),
    .INIT_10(256'hFFFF37657CD5C06881DABCBEAD555555555555555554655555555C37FFFFFF53),
    .INIT_11(256'hFFFF4F589CD5C17DF2D8BDCFA75555555555555555D99D55555555B7FFFFFFD4),
    .INIT_12(256'hFFFFD5F1ACD5C3FFD6FA8BD09B555555555555555746D555555555B7FFFFFFF4),
    .INIT_13(256'hFFFFF9DF64D5E3FFF6D002FFA6D55555555555555F1B555555555507FFFFFFFD),
    .INIT_14(256'hFFFFF569FAD5EBFFF65AF827CA75555555555555784555555555572FFFFFFFFF),
    .INIT_15(256'hFFFFFDE8F0D5E3FFF668F580F335545555555555E93D7FFF5555556FFFFFFFFF),
    .INIT_16(256'hFFFFFF66D6D5EBFFFE66FF681E6D54D55555555796AAA80F55F55567FFFFFFFF),
    .INIT_17(256'hFFFFFF66DC55EBFFFCCDFFF60DE75FD55555555C580F555557F55547DD5FFFFF),
    .INIT_18(256'hFFFFFFE43E55E7FFFD4FFFDF68935955515555D1AFF57D5FFD6555CF9F7FFFFF),
    .INIT_19(256'hFFFFFFFF9EF5E7FFFFAFFD17FE36D155FB55574D9200000027D555C592DFFFFF),
    .INIT_1A(256'hFFFFFFEF2FB5C7FFFD1FFD7DFE0C5355C5555D328008280802BD55E58E1FFFFF),
    .INIT_1B(256'hFFFFFFFDAD35C7FFFFBFFEF7FD0F135545555660009FFFFF682755E91DBFFFFF),
    .INIT_1C(256'hFFFFFFDCC335CBFFFFBFF6FDFF0B8F554D55F7887557FFFFDD0355E6B73FFFFF),
    .INIT_1D(256'hFFFFFFD5FBB5E3FFFF1FF77DFFEAC755CD57B4155FFFFFFD7F07556E5617FFFF),
    .INIT_1E(256'hFFFFFFD47A35F3FFFFBFF777FFE86F55ED76E17E67FFFFFFFC2D556E7297FFFF),
    .INIT_1F(256'hFFFFFFE47C155BFFFF7FF657FFC22757ADDB25F6F7FFFFFFF43D55FEDBD7FFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n653,addra[14:13]}),
    .dia({open_n657,open_n658,open_n659,open_n660,open_n661,open_n662,open_n663,1'b0,open_n664}),
    .rsta(rsta),
    .doa({open_n679,open_n680,open_n681,open_n682,open_n683,open_n684,open_n685,open_n686,inst_doa_i1_002}));
  // address_offset=8192;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hBBCEEAF85003914557AB6C85555555555555555555A441214A84040000000000),
    .INIT_01(256'hFBBD0AB90403E15557EB6C95555555555555555554357DB553AC050000000000),
    .INIT_02(256'hAAFBFBBF4400D1555728198555555555555555555520B18554B0000000000034),
    .INIT_03(256'h2AFBBA7E440F1555532D0E15555555555555555555491655552F000000000265),
    .INIT_04(256'h7FFFBFCF4573255552681E51555555555555555555560B155537C00000000035),
    .INIT_05(256'hFBFBBFCA140B9555537C96115555555555555555154749555143B000000000EA),
    .INIT_06(256'hEEB0FE9294F4555557F9D655555555555555555555529915551AEC000000008C),
    .INIT_07(256'hF5BA7AF6D625555542E4AB1555555555555555555555DD515112A7000143C400),
    .INIT_08(256'hFE3CCEE4C531555552A188C55555555555555555555591145D44F4000000CC40),
    .INIT_09(256'hFEEE3BA14621555552B0961555555555555555555555854226E4C300000029C0),
    .INIT_0A(256'hFF6A8AF95291504157E1CAB155555555555555555554D05DD5481300005183CA),
    .INIT_0B(256'hFFF2C8F9D1C505A847F63DFD15555555555555555554003645143380000B2B79),
    .INIT_0C(256'hFFEBDB7C5E85411AACFE606D54555555555555555550568D5555437000050FF1),
    .INIT_0D(256'hFFF0ABCE4D9544001C37712F555555555555555555555BA555555B60000533FE),
    .INIT_0E(256'hFFFBE7324FC53B540A22F40E84555555555555555550638555554904000504BF),
    .INIT_0F(256'hFFFDBD8146552005386BEC17C5555555555555555554FA55555441B40005432B),
    .INIT_10(256'hFFFF897FC755727A503EDB83E555555555555555554674555554534D000055DF),
    .INIT_11(256'hFFFFFDDAB30531974A32D5F9E055555555555555151485555555555800004533),
    .INIT_12(256'hFFFFC6193605304022135D4FD855555555555555146255555555554800000048),
    .INIT_13(256'hFFFFFA4C121503EFFA5E80971715555555555555529855555555546800000002),
    .INIT_14(256'hFFFFF8E9771507FFF9C900007B055515555555554B3005555555548000000000),
    .INIT_15(256'hFFFFFD3B0E111BFFFCAEBC035DC55755555555552DC155555555547440000005),
    .INIT_16(256'hFFFFFE2400411BFFF9A6FFF04261521555555554C09017EE1105546C11400000),
    .INIT_17(256'hFFFFFFC1C3140FFFFA65FFFE5D354E155155505652FF505152B5552822F00000),
    .INIT_18(256'hFFFFFFF2820403FFFD7BFFBBB6F849155855541CB100694151615530F4900000),
    .INIT_19(256'hFFFFFFFB16C507FFFDAFFFC3E1521D552C555470D8100001A5455521AD200000),
    .INIT_1A(256'hFFFFFFEEE38537FFFECFFD26FE6B5D557515509C4006EBA501945125EEF50000),
    .INIT_1B(256'hFFFFFFEA808133FFFE0FFE39FE10C855205546D0068155556401553814000000),
    .INIT_1C(256'hFFFFFFDEA9952FFFFE5FFE6CBF82E855255525065EB950042508552794900000),
    .INIT_1D(256'hFFFFFFD2B7857FFFFFFFFE2DFF07C154F141959BFFFFFAAF8541553707D80000),
    .INIT_1E(256'hFFFFFFC2B8D57BFFFFAFFB5AFF9DB854B1566DAA7FFFFFFFF50055365E980000),
    .INIT_1F(256'hFFFFFFF2BB5153FFFFEFFB46BFFAF054F159BEB7B3FFFFFFFF21557655880000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n712,addra[14:13]}),
    .dia({open_n716,open_n717,open_n718,open_n719,open_n720,open_n721,open_n722,1'b0,open_n723}),
    .rsta(rsta),
    .doa({open_n738,open_n739,open_n740,open_n741,open_n742,open_n743,open_n744,open_n745,inst_doa_i1_003}));
  // address_offset=8192;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hAE162AABAFFF4FEFFC7AAB3FFFFFFFFFFFFFFFFFFF16A3DFE0ABFBFFFFFFFFFF),
    .INIT_01(256'hAAE13FABFBFF1BFFFD7BAE3FFFFFFFFFFFFFFFFFFEDCD64FF86FFAFFFFFFFFFF),
    .INIT_02(256'hEAAE4FAABBFE3FFFFCFBFE6FFFFFFFFFFFFFFFFFFF8B0B2FFE5FFFFFFFFFFFFF),
    .INIT_03(256'hFAAAFAFBBBFCFFFFF9BEFDFFFFFFFFFFFFFFFFFFFFF2BCBFFFC7FFFFFFFFFFCA),
    .INIT_04(256'hAAAAAABBBABCDFFFF9BFFCFFFFFFFFFFFFFFFFFFFFF8A1BFFF80FFFFFFFFFFC6),
    .INIT_05(256'h9AAEAAFEEBF57FFFF8EB69BFFFFFFFFFFFFFFFFFFFFDB3FFFBE43FFFFFFFFFE4),
    .INIT_06(256'hF7ABAABEABC1FFFFFDAB79BFFFFFFFFFFFFFFFFFFFF933FFFFF15FFFFFFFFFFF),
    .INIT_07(256'hFAECEAAAAB82FFFFEDEF71BFFFFFFFFFFFFFFFFFFFFE33FFFBF91BFFFEBFFBFF),
    .INIT_08(256'hFDEA6ABBFADFFFFFF9AE726FFFFFFFFFFFFFFFFFFFFF2BBEF2EE5BFFFFFD7FBF),
    .INIT_09(256'hFE2BDEAEBBCBFFFFFCFE21ABFFFFFFFFFFFFFFFFFFFF6FE88D1E0BFFFFFD06FF),
    .INIT_0A(256'hFFCEE7AAAF3BFFEBF8FE204FFFFFFFFFFFFFFFFFFFFE3FE33FE787FFFFAE392B),
    .INIT_0B(256'hFFDFB6EEAF2FFF13A9ED9256FFFFFFFFFFFFFFFFFFFFFE8CEFFF90BFFFFF8F97),
    .INIT_0C(256'hFFE2A1FBAD2FFFE447ED9E87FFFFFFFFFFFFFFFFFFFFF973FFFFF1BFFFFAE2F9),
    .INIT_0D(256'hFFFFE56EBD6FEAAAB7E98B95FFFFFFFFFFFFFFFFFFFFF10FFFFFF4FFFFFAF8BF),
    .INIT_0E(256'hFFFDECDEBC2F91BBB0BC5AF46EFFFFFFFFFFFFFFFFFAC92FFFFFE0FBFFFAFE7F),
    .INIT_0F(256'hFFFE7A7EBCBF900142F503BD6FFFFFFFFFFFFFFFFFFF44FFFFFFE87BFFFABF8B),
    .INIT_10(256'hFFFF2BDFF9FFD09002E175780FFFFFFFFFFFFFFFFFE99AFFFFFFF97AFFFFAAF6),
    .INIT_11(256'hFFFF9BF479AF92BFF1E12B434AFFFFFFFFFFFFFFFFB72BFFFFFFFF2FFFFFBAF9),
    .INIT_12(256'hFFFFFFF658AF92FFEDF453B467FFFFFFFFFFFFFFFE98BFFFFFFFFF7FFFFFFFBA),
    .INIT_13(256'hFFFFF6E7C9BF96FFF9F551284DBFFFFFFFFFFFFFF837FFFFFFFFFF1BFFFFFFFE),
    .INIT_14(256'hFFFFFE9695BF93FFFDA5E00FC5EFFEFFFFFFFFFFE48EAFFFFFFFFE4FFFFFFFFF),
    .INIT_15(256'hFFFFFF90A5BF83FFFDD5EA00E63FFDFFFFFFFFFF872BFFFFFFFFFE9BBFFFFFFA),
    .INIT_16(256'hFFFFFF9DE9FF83FFF989FE902CCBF9BFFFFFFFFE7C040455AFAFFEDFEEBFFFFF),
    .INIT_17(256'hFFFFFF8868BF97FFFD9BFFF943CFE0BFFFFFFFFDE144EFFEA90FFFCEFFAFFFFF),
    .INIT_18(256'hFFFFFFD968EF9BFFFF9AFFFF9122E7BFE6FFFFA21ABB82AFAB8FFF8B3FEFFFFF),
    .INIT_19(256'hFFFFFFC1696F9BFFFF4FFE2FED3DB6FF86FFFEDE255000044FAFFF9E24BFFFFF),
    .INIT_1A(256'hFFFFFFC45C6F9BFFFF6FFEBAF90DA7FFDFFFFB3500044140017FFF8E043AFFFF),
    .INIT_1B(256'hFFFFFFC44E2F8BFFFE6FFDBBFF4A22FFDFFFE890047FFFFE801BFF862A3FFFFF),
    .INIT_1C(256'hFFFFFFE0137F97FFFF3FF9FFFF5342FF9FFF8F01EBEBFFFBEF42FF982E7FFFFF),
    .INIT_1D(256'hFFFFFFFC113FC3FFFF3FFDAEBF958FFE1BEB6D7AFFFFFFFBBE1BFF8DE92FFFFF),
    .INIT_1E(256'hFFFFFFFC152FC7FFFF2FFCA8BF80C6FE0BE883ADCBFFFFFFEF1BFF88E52FFFFF),
    .INIT_1F(256'hFFFFFFDC106BE2FFFFBFFCBCFFD11EFE4BF30FF8BBFFFFFFFC0BFFC8A76FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n771,addra[14:13]}),
    .dia({open_n775,open_n776,open_n777,open_n778,open_n779,open_n780,open_n781,1'b0,open_n782}),
    .rsta(rsta),
    .doa({open_n797,open_n798,open_n799,open_n800,open_n801,open_n802,open_n803,open_n804,inst_doa_i1_004}));
  // address_offset=8192;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h565D7F7DFFFF721AA15C6B2AAAAAAAAAAAAAAAAAA02C4B909B89FFFFFFFFFFFF),
    .INIT_01(256'hF56DB6FDF5FD46AAA2DD4F2AAAAAAAAAAAAAAAAAA95E09BAAE8FF7FFFFFFFFFF),
    .INIT_02(256'h7FDC1E9C7DFD4AAAAA15DC3AAAAAAAAAAAAAAAAAA86E9712AB277FFFFFFFFF5F),
    .INIT_03(256'h7FFD6DEC57DFCAAAA57B7DEAAAAAAAAAAAAAAAAAAAACE002AA337FFFFFFFFF70),
    .INIT_04(256'hAFFDFD947FD052AAA7DB2DAAAAAAAAAAAAAAAAAAAAA4FC6AAA507FFFFFFFFFE8),
    .INIT_05(256'hDDF3F79B7F5DEAAAAD7345EAAAAAAAAAAAAAAAAAAAA380AAAE0E7FFFFFFFFF47),
    .INIT_06(256'hEFDF7FDD9F548AAA8013A062AAAAAAAAAAAAAAAAAAA676AAAAA457FFFFDFFDFE),
    .INIT_07(256'h767377469DDA2AAAB2B51E6AAAAAAAAAAAAAAAAAAAA1B6A00C845BFFFF7DDFFD),
    .INIT_08(256'h7DFC0FCF5F7EAAA2A85D185AAAAAAAAAAAAAAAAAAAA100C8FC117FFFFFDBF77F),
    .INIT_09(256'hFF77A9F75F0EAAA285CFFC1CAAAAAAAAAAAAAAAAAAA15AB96DFB0FFFFFF53DFF),
    .INIT_0A(256'hFF472659FFD6AA3C8744C20AAAAAAAAAAAAAAAAAAAA02A14088C17FFFFF71EFB),
    .INIT_0B(256'hFDFD66397C1AA10DB767A7932AAAAAAAAAAAAAAAAAAA81D01A0073BFFFFDCB62),
    .INIT_0C(256'hFFD55F25F55AA225A0ECAB372AAAAAAAAAAAAAAAAAAA8662AAAAA93FFFFFF2DD),
    .INIT_0D(256'hFFF2DFD85DDA35FF64ED9C4D2AAAAAAAAAAAAAAAAAAA038AAAAA821FFFFFFC3D),
    .INIT_0E(256'hFFF69D9CFD5AC87A7E805D0493AAAAAAAAAAAAAAAA85999AAAAA9E7FFFFFFD2F),
    .INIT_0F(256'hFFFDD17FF72A600076865245C0AAAAAAAAAAAAAAAA80842AAAAA985FFFFFFFF7),
    .INIT_10(256'hFFFF45B5760A0034E04D458C8AAAAAAAAAAAAAAAAABA37AAAAAAAE17FFFFFFC3),
    .INIT_11(256'hFFFF85DFF4DA629F7D4846BCC5AAAAAAAAAAAAAAAA580CAAAAAAA9F7FFFFFFDA),
    .INIT_12(256'hFFFFCA422DDA41FFC15F80EF442AAAAAAAAAAAAAA16CA2AAAAAAA8C5FFFFFDFA),
    .INIT_13(256'hFFFF5E63BB4A69755162237F9BCAAAAAAAAAAAAAAD660AAAAAAAAAE1FFFFFFFC),
    .INIT_14(256'h557FF0B8E56A4FFFF3ADF80D1572A82AAAAAAAA83B5178AAAAAAA9DFFFFFFFFF),
    .INIT_15(256'hFFFFFE79DA6A6BFFF31E50C19FEAAA2AAAAAAAAA445CA8AA0AA2AB7FFFFFFFFD),
    .INIT_16(256'hFFFFFD13B8226FFFFD93FFB46806A0CAAAAAAA8BC8B801412AFAAB777FFFFFFF),
    .INIT_17(256'hFFFFFFAA972A67FFF46EF7F1007E1FEAAAAAAA2BA361EAA88B7AAAB75FFFFFFF),
    .INIT_18(256'hFFFFFFF31EFA4BFFFE0DF7B5BC6D396A83AAA8C7976BF5E054B2AA54F7FFFFFF),
    .INIT_19(256'hFFFFFDC0CE1A6BFFFFFFFEA3D71846AAFB2AA34E3C4000092CFAAA7A4B7FFFFF),
    .INIT_1A(256'hFFFFFFCD271A63FFFE0FFFF4FD860CAA9C2AAF71C02A16A6038AAAC47A3FFFFF),
    .INIT_1B(256'hFFFFFFCDBA1A7BFFFF7FF834FE2C41AA3AAA3CB022657FF79C34AACCFE9FFFFF),
    .INIT_1C(256'hFFFFFFCFDE62D7FFFF5FF2FC7F8F5DA81AAA5B445A2B5FDDE4078AC31927FFFF),
    .INIT_1D(256'hFFFFFFE54800A7FFFF8FF4FEFFF5FEA976B4902A4FFFDFD4B780AA439247FFFF),
    .INIT_1E(256'hFFFFFFCF604A1BFFFFFFFC817FF31FA94432D29253FFFFFFF72EAAEE9EA7FFFF),
    .INIT_1F(256'hFFFFFFF74C6629FFFF1FF6817FC8FFAB24211E7CEBFFFFFFF81EA88C7C0FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n830,addra[14:13]}),
    .dia({open_n834,open_n835,open_n836,open_n837,open_n838,open_n839,open_n840,1'b0,open_n841}),
    .rsta(rsta),
    .doa({open_n856,open_n857,open_n858,open_n859,open_n860,open_n861,open_n862,open_n863,inst_doa_i1_005}));
  // address_offset=8192;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h77CDD7D600024F555CD71C9555555555555555555789FEF75BE2000000000000),
    .INIT_01(256'h5776E5D40A00C5555ED4123555555555555555555711B32D5478080000000000),
    .INIT_02(256'h5577F7770202D5555E1628355555555555555555556B8E1D551A80000000008A),
    .INIT_03(256'h355777BD28291555571C8BB55555555555555555555D7CFD55D6800000000252),
    .INIT_04(256'h1D5757EF00000D555794AB555555555555555555557270555579000000000038),
    .INIT_05(256'hFF5555CD80AF55555FBEC9D555555555555555555557D35555DBC00000000095),
    .INIT_06(256'hF770D5614019F5555FF6485D55555555555555555556A3555573F00000200008),
    .INIT_07(256'hF855B5F1C295D55555DAE7555555555555555555555E2B57FF54720000002002),
    .INIT_08(256'hFD3DDD70209B55555F50E4555555555555555555555C975F0BF5D8000020C000),
    .INIT_09(256'hFDFF3F582205555573F0612D5555555555555555555CD577282F3200000A5400),
    .INIT_0A(256'hFF8545F402CD55FF71D840455555555555555555555DB5643F596800000AC3E6),
    .INIT_0B(256'hFFF1C4F480155E02F9F931795555555555555555555555B2F57D73400002173E),
    .INIT_0C(256'hFFD747BE0155555A04FB3574D555555555555555555556EB55555C2000008FF2),
    .INIT_0D(256'hFFF057CF2AD575FFDC38954D55555555555555555555D18D55557F20000023FD),
    .INIT_0E(256'hFFF7FB330B35C82D7A11DF7E15555555555555555557F395555556800000087F),
    .INIT_0F(256'hFFFC7E400BD55000BC97DB71DD55555555555555555FC655555574400000021F),
    .INIT_10(256'hFFFF56B009D55397023753BE8555555555555555557F9355555557A8000000AF),
    .INIT_11(256'hFFFFF69F41D5726AAD3DDF196155555555555555554CBD5555555C2800000001),
    .INIT_12(256'hFFFFC90FFBD57080112389FF6FD555555555555555BA75555555572800000206),
    .INIT_13(256'hFFFFF58B415553DFF5ADC09C695555555555555556EDF5555555559400000001),
    .INIT_14(256'hFFFFF4FB4B555BFFF6C60C3977B5575555555555599F5555555555C000000000),
    .INIT_15(256'hFFFFFE335D5577FFFC5D7C03DCF554D555555555467757FFF555571800000000),
    .INIT_16(256'hFFFFFD3275DD77FFF659FDD03E8D54D555555557EB3575405DF5553080000000),
    .INIT_17(256'hFFFFFFF715557FFFF59AFFF7A01378D55D55555D8F60355F5E25555A20000000),
    .INIT_18(256'hFFFFFFD5FE3553FFFEB7FF6F53D572D5735555DEB7FE281DF765557AC8800000),
    .INIT_19(256'hFFFFFFCC1E155BFFFE5FFD6BD02A7755CB555738A5000008C175555056A00000),
    .INIT_1A(256'hFFFFFFE24E957BFFFDCFFDFBFD175F55DB555EEC0009D75A029D55C4F8400000),
    .INIT_1B(256'hFFFFFFC0BD9553FFFD0FFF36FF01F955555572E00142AAAA982355E687E00000),
    .INIT_1C(256'hFFFFFFE237F5DFFFFDAFFFF4FFC151577D554A096576A0083A8555E315C80000),
    .INIT_1D(256'hFFFFFFC82435C7FFFFFFF9DEFFA1E357155F8847BFFFF55F60AF5569D6680000),
    .INIT_1E(256'hFFFFFFCA0BD5C7FFFF5FF16D7F427357057C96577FFFFFFFDB1555E05C880000),
    .INIT_1F(256'hFFFFFFD2003DF7FFFFDFF3DDFFD85357876A79F55BFFFFFFFF2D55C0CB080000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n889,addra[14:13]}),
    .dia({open_n893,open_n894,open_n895,open_n896,open_n897,open_n898,open_n899,1'b0,open_n900}),
    .rsta(rsta),
    .doa({open_n915,open_n916,open_n917,open_n918,open_n919,open_n920,open_n921,open_n922,inst_doa_i1_006}));
  // address_offset=8192;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5D291757FFFF8FFFFF35D7FFFFFFFFFFFFFFFFFFFF5151EFD65FFFFFFFFFFFFF),
    .INIT_01(256'h55D29FD5FFFD17FFFDB5D5FFFFFFFFFFFFFFFFFFFFC645DFF79FFFFFFFFFFFFF),
    .INIT_02(256'hD55D8F55FFFD1FFFFFF7FF7FFFFFFFFFFFFFFFFFFF57775FFD6FFFFFFFFFFFDF),
    .INIT_03(256'hD555F5F7FFFC5FFFF47FFCFFFFFFFFFFFFFFFFFFFFF37D7FFFE3FFFFFFFFFF0D),
    .INIT_04(256'h55555577FFDD7FFFF67FFEFFFFFFFFFFFFFFFFFFFFFD757FFF627FFFFFFFFFCB),
    .INIT_05(256'h6D5D55F5FFF0BFFFFED7B4FFFFFFFFFFFFFFFFFFFFF677FFFFF01FFFFFFFFFD8),
    .INIT_06(256'hD957557D7F60FFFFFC57157FFFFFFFFFFFFFFFFFFFF777FFFFFCA7FFFFFFFFFF),
    .INIT_07(256'hF5DCD55D7F43FFFFFCDFB07FFFFFFFFFFFFFFFFFFFFFF7FFFFF52FFFFFFD7FFF),
    .INIT_08(256'hFED5957F7FEFFFFFF45FB19FFFFFFFFFFFFFFFFFFFFD77FD55FD27FFFFFEB7FF),
    .INIT_09(256'hFD35E55FFFF7FFFFF67D127FFFFFFFFFFFFFFFFFFFFD9FF6DF57E7FFFFFE0B7F),
    .INIT_0A(256'hFFDDDB57FF9FFFFFFCFF9F9FFFFFFFFFFFFFFFFFFFFD7F73FFD769FFFFFD3617),
    .INIT_0B(256'hFFEF79DFFD5FFF777EDE6DA5FFFFFFFFFFFFFFFFFFFFFD4FFFFF407FFFFF4FEB),
    .INIT_0C(256'hFFD1F2F7F69FFFDDDBDECFE9FFFFFFFFFFFFFFFFFFFFF71FFFFFF8FFFFFFD1F6),
    .INIT_0D(256'hFFFFDA9DFE9FF5FFF3D447527FFFFFFFFFFFFFFFFFFFDEFFFFFFF07FFFFFF47F),
    .INIT_0E(256'hFFFEDCEDFCFFD5F7577CA7F35FFFFFFFFFFFFFFFFFFFE65FFFFFD8FFFFFFFDBF),
    .INIT_0F(256'hFFFFB5BFFE7F400229FA25763FFFFFFFFFFFFFFFFFFF1B7FFFFFF49FFFFFFF47),
    .INIT_10(256'hFFFF17E576FF606001D09EF7F7FFFFFFFFFFFFFFFFF46FFFFFFFF4BFFFFFFFF9),
    .INIT_11(256'hFFFF6FC296FF417FDADA3765BDFFFFFFFFFFFFFFFF53DFFFFFFFFD1FFFFFFFD6),
    .INIT_12(256'hFFFFFFD126FF41FFDEF8AD5A93FFFFFFFFFFFFFFFDCFFFFFFFFFFFBFFFFFFFF7),
    .INIT_13(256'hFFFFF9D5C47F49FFF6FAA0570E7FFFFFFFFFFFFFF5B3FFFFFFFFFFA7FFFFFFFD),
    .INIT_14(256'hFFFFFD4D587F43FFFE5AD82F6AFFFDFFFFFFFFFFDCCFFFFFFFFFFD8FFFFFFFFF),
    .INIT_15(256'hFFFFFF4E507F63FFFEEAD502F1BFFFFFFFFFFFFF7B17FFFFFFFFFFE7FFFFFFFF),
    .INIT_16(256'hFFFFFF4CF4FF63FFF646FF601FF7F7FFFFFFFFFF16CAA23757FFFF47FFFFFFFF),
    .INIT_17(256'hFFFFFF64567F6BFFFE67FFFE87C7F5FFF7FFFFFCDA175FF55D5FFFEDFFFFFFFF),
    .INIT_18(256'hFFFFFFE61DFF47FFFF65FF5F6019FFFFDFFFFFFBCD77D7DD577FFF671FFFFFFF),
    .INIT_19(256'hFFFFFFDDBF5F47FFFF8FFF3FDEB771FFDFFFFF45F0200000357FFF4F187FFFFF),
    .INIT_1A(256'hFFFFFFFDB5DF47FFFF9FFC35F60CFBFFCFFFFFBA0008828000DFFFF3279FFFFF),
    .INIT_1B(256'hFFFFFFDDED5F67FFFD9FF6F5FD8595FFEFFFFF6000BFFFFD400FFFF9B5BFFFFF),
    .INIT_1C(256'hFFFFFFDF6BBFCBFFFF3FFE3DFF23A5FF6FFF570217D7FFF7FF89FFFCDD1FFFFF),
    .INIT_1D(256'hFFFFFFFD59FFF3FFFF3FF4BF7FCA6FFFC7FFDCB77FFFFFF75D07FF7E7F3FFFFF),
    .INIT_1E(256'hFFFFFFFF5EBFF3FFFF1FF4BCFF4ECFFF77F76B54A7FFFFFFDE07FFF7D3FFFFFF),
    .INIT_1F(256'hFFFFFFE7571FD9FFFF7FF6A0FFEF2FFFF75F0FF2D7FFFFFFFC1FFFD7737FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_008192_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n948,addra[14:13]}),
    .dia({open_n952,open_n953,open_n954,open_n955,open_n956,open_n957,open_n958,1'b0,open_n959}),
    .rsta(rsta),
    .doa({open_n974,open_n975,open_n976,open_n977,open_n978,open_n979,open_n980,open_n981,inst_doa_i1_007}));
  // address_offset=16384;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFD0C42D59DFFFFFF100FFE0C3DDFB4E8FDD7FFFFFFFFD17F5C9C027FFFF),
    .INIT_01(256'hFFFFFFC6D689D7DFFFFFF906FFC42355B5E53FFFF3FFFFFFF807F5E0B387FFFF),
    .INIT_02(256'hFFFFFFCCE291FCFFFFFFFD677FF681B87719FFD477FFFFFFF837FD54CD37FFFF),
    .INIT_03(256'hFFFFFFFC6159FB3FFFFFFF3D7FEE5D4ED26BFFE219FFFFFFF3D7FD39BD37FFFF),
    .INIT_04(256'hFFFFFFF19A597F8FFFFFFFFFFFFF9EF16EBFFFF00BFFFFFFD937FF9E39D15FFF),
    .INIT_05(256'hFFFFFFFB1A8F7753FFFFFFFFFDB5B7D0F993FFD027FFFFFFFB5FFF2A1FF09755),
    .INIT_06(256'hFFFFFFFDA76755DCFFFFFFFFF6F57DFDD8EFFFE83BFFFFFFEC57FD3A0CC509F0),
    .INIT_07(256'hFFFFFFFF0C77557D7FFFFFFF6BF5FFF571FFFFD8B7FFFFFF175FDC84AA0765C0),
    .INIT_08(256'hFFFFFFFF2881555D7BFFFFFDAFFFFFFD7F6FDFF7AFFFFFFFA55DD13BB6BB47FF),
    .INIT_09(256'hFFFFFFFF8FEE5557491FFF0CDDFFFFFDFD6FFFFCBFFFFFFDFD5FD7ABB6C7C7FF),
    .INIT_0A(256'hFFFFFFFFF3E65555768E3707557FF7FD7DCFFFFFFFFFFFFFBD5F755046BBF67F),
    .INIT_0B(256'hFFFFFFFFD286555555582DD5557FFDFD7DD9FFFFFFFFFFFD7FD75032E715167F),
    .INIT_0C(256'hFFFFFFFFFEB9555FFFFFFD57F57FFF7D7D77FFFFFFFFFFF03FF75F10EB8B9DBF),
    .INIT_0D(256'hFFFFFFFFFFD3FFFFFFFFFD7FFFFFF7F7FFFD7FFFFFFFFFE3FFFDFF717753DDBF),
    .INIT_0E(256'hFFFFFFFFFF04FFFFFFFFFFFFFFFFDAD7FFF747FFFFFFFFF9FFF5351332F547BF),
    .INIT_0F(256'hFFFFFFFFFF4EFFFFFFFFFFFFFFFF6ED7FFF5DBFFFFFFFF1D7FF7792E88F7355D),
    .INIT_10(256'hFFFFFFFFFF711FFFFFFFFFFFFFFF245FFFF574BFFFFFFEBD7FD5A7B0F3FF9F97),
    .INIT_11(256'hFFFFFFFFF1B99FFFFFFFFFFFFFFFA47FFFFDDD0BFFFFCD77FFFE42034FF72F8F),
    .INIT_12(256'hFFFFFFFF6F9A97FFFFFFFFF555F76ED7FFFFF72CA9ACE9F7FFDE0EC49FFFDFE2),
    .INIT_13(256'hFFFFFFFFCA60D5FFFFFFFFF555F7E1FFFFFFF5DF882447FFFFDE73A2FFFF7373),
    .INIT_14(256'hFFFFFFCD0B89B5FFFFFFFFFFFFFFF7FD555555FD7DD757FFFFD47E9D3FFFD0DF),
    .INIT_15(256'hFFFFFF946F15057FFFFFFFF55557FD041D757575555557FFFF553053A257F57D),
    .INIT_16(256'hFFFFFFFFFCE2E57FFFFFFFD57F05D2F68172D9F5FFFFFFFFFD57C9FA80E5F637),
    .INIT_17(256'hFFFFFFFFF44A357FFFFFFF41C389C169AFF410B5FFFFD7FFFDF737FFFF975FED),
    .INIT_18(256'hFFFFFFFF80B7DD7FFFFF5CD3C9385FFFFFFFFB6DFFFF57FFF56579FFFFDB84D7),
    .INIT_19(256'hFFFFFFDF5E8FA57FFFDD0346FFFFFFFFFFFFFF27FFFFFFFFD6912CFFFFFD2567),
    .INIT_1A(256'hFFFFFD4D6EFB717FFFD5C3FFFFFFFFFFFFFFFFA2D5FFFFFFD771AC7FFFFFF4DD),
    .INIT_1B(256'h0AA06A254AEA6F7FFFD5D3FFFFFFFFFFFFFFFFB1B5FFFFFF51D643FFFFFFFFFF),
    .INIT_1C(256'h00C2B16AA88AF85FFF55C5E4FFDC377588BCFFB765FFFFFF7BD51C7FFFFFFFFF),
    .INIT_1D(256'h55556AAA8AA95EDFFFD64F1AAAAAAAEAAAA55B99397FFFFD52B5764FFFFFFFFF),
    .INIT_1E(256'hAAAAAAAAAAA9FA57FDF4E67FD55555555575679D7D5FFFFD5C54133DFFFFFFFF),
    .INIT_1F(256'hAAAAAAAAAAA15C97FDF41FFD5D5577FF5295DD77C65FFFDFEBC8B30FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1007,addra[14:13]}),
    .dia({open_n1011,open_n1012,open_n1013,open_n1014,open_n1015,open_n1016,open_n1017,1'b0,open_n1018}),
    .rsta(rsta),
    .doa({open_n1033,open_n1034,open_n1035,open_n1036,open_n1037,open_n1038,open_n1039,open_n1040,inst_doa_i2_000}));
  // address_offset=16384;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFD0C64A8EFFFFFFF7A2FFEC72885E6277DEF1FFFFFFF48AAA8B2782AAAA),
    .INIT_01(256'hFFFFFFCCD46E8DFFFFFFFDADFFF69B18BDA8FFE6F5FFFFFFF4DAAA88C682AAAA),
    .INIT_02(256'hFFFFFFDEC0D6A97FFFFFFEEBFFF00B7982F4FFCEF9FFFFFFF8AAAA85A232AAAA),
    .INIT_03(256'hFFFFFFFE4196A7BFFFFFFF5FFFDA6B2D91C7FFE053FFFFFFFE2AAA041A32AAAA),
    .INIT_04(256'hFFFFFFF91176AA7FFFFFFFFFFF4828A6061BFFE283FFFFFFF94AAA883A360AAA),
    .INIT_05(256'hFFFFFFFF9312AABFFFFFFFFFFFEAAA80A19FFFC2A3FFFFFFC2AAAA8C3A14CA00),
    .INIT_06(256'hFFFFFFFF2412AAADFFFFFFFFFFAAAAAAA2BFFFFA97FFFFFFDDAAAA141130D3F2),
    .INIT_07(256'hFFFFFFFE6E3AAAA93FFFFFFFF2AAAAAAA2BFFFDA9FFFFFFFE2AAA8143532B77F),
    .INIT_08(256'hFFFFFFFFE220AAA857FFFFF4AAAAAAAAAA9FFFF9DFFFFFFFA2A8A703059627FF),
    .INIT_09(256'hFFFFFFFFDAC5AAAA077FFFE68AAAAAAAAABFFFFFFFFFFFFDCAAAA1F3094294FF),
    .INIT_0A(256'hFFFFFFFFD185AAAAA25EA282AAAAAAAAAA83FFFFFFFFFFFE8AAAA99051C6AB7F),
    .INIT_0B(256'hFFFFFFFFDF8DAAAAA82AA2AAAAAAAAAAAAA6FFFFFFFFFFF72AAA8992426E60FF),
    .INIT_0C(256'hFFFFFFFFF064AAAAAAAAAAAAAAAAAAAAAAA3BFFFFFFFFFF26AAA8C7047D708EF),
    .INIT_0D(256'hFFFFFFFFFD8EAAAAAAAAAAAAAAAAA8AAAAA8EFFFFFFFFFDCAAAAA2F14A80389F),
    .INIT_0E(256'hFFFFFFFFFCBCAAAAAAAAAAAAAAAAA2AAAAAA3BFFFFFFFFF0AAAA535386A9FC53),
    .INIT_0F(256'hFFFFFFFFFDF6AAAAAAAAAAAAAAAA8CAAAAAA84FFFFFFFF12AAAA04CC79A3B72F),
    .INIT_10(256'hFFFFFFFFFD196AAAAAAAAAAAAAAA8C2AAAAAA13FFFFFFC4AAAA8833BD6AADDCC),
    .INIT_11(256'hFFFFFFFFFD8D6AAAAAAAAAAAAAAA0E2AAAAAA8F7FFFFDF2AAAA9B80F5AAA8FD9),
    .INIT_12(256'hFFFFFFFFEE456AAAAAAAAAAAAAAA06AAAAAAAAE39DD0D8AAAAAAEC3F4AAABFF6),
    .INIT_13(256'hFFFFFFFC438FAAAAAAAAAAAAAAAAA2AAAAAAAA895D5E92AAAAA97A55AAAA0BFA),
    .INIT_14(256'hFFFFFF60DEE52AAAAAAAAAAAAAAAAAAAAAAAAAA82A82AAAAAAA869C46AAA81FD),
    .INIT_15(256'hFFFFFFF43D619AAAAAAAAAAAAAAAA8514AA02AAAAAAAAAAAAAAA2544E7AAABFF),
    .INIT_16(256'hFFFFFFFFFEF4DAAAAAAAAAAAAA50A27D7F7D64AAAAAAAAAAAAAA97FD3EBAA03F),
    .INIT_17(256'hFFFFFFFFF713CAAAAAAAAA148B5E9DCA77F59C6AAAAAAAAAAAAA7BFFF9F20AFF),
    .INIT_18(256'hFFFFFFFFE55D6AAAAAAA08769F8F7FFFFFFFF55AAAAAAAAAA89885FFFF630997),
    .INIT_19(256'hFFFFFFF96EE522AAAAA897E97FFFFFFFFFFFFF12AAAAAAAAA9546EFFFFFF6DD7),
    .INIT_1A(256'hFFFFF6F65B9D3EAAAAA847FFFFFFFFFFFFFFFFEDAAAAAAAAAA8D93FFFFFFFD83),
    .INIT_1B(256'hAAAAF795477F92AAAAA8C7FFFFFFFFFFFFFFFFC16AAAAAAAA5CC253FFFFFFFFF),
    .INIT_1C(256'h00C0AD7FDDDD99AAAAA849D0557C8A28A28B7FC8DAAAAAAAA6B040FFFFFFFFFF),
    .INIT_1D(256'h55557FFFDFFC8DAAAAA9E9CAAAAAAAAAAAA09F6C96AAAAAA836035BFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFE2C2AAAA962000000000000002A7828AAAAAA8D066E7FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFEA36AAAA94000280022AA054208402DAAAAAAABFDCA17FFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1066,addra[14:13]}),
    .dia({open_n1070,open_n1071,open_n1072,open_n1073,open_n1074,open_n1075,open_n1076,1'b0,open_n1077}),
    .rsta(rsta),
    .doa({open_n1092,open_n1093,open_n1094,open_n1095,open_n1096,open_n1097,open_n1098,open_n1099,inst_doa_i2_001}));
  // address_offset=16384;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFE73B157BFFFFFFF655FFD9A557AD9C1FF1FFFFFFFFFE355556C3D7FFFF),
    .INIT_01(256'hFFFFFFDB2B357AFFFFFFF659FFDBCCE7CAFA7FF9F7FFFFFFF4355555A1D7FFFF),
    .INIT_02(256'hFFFFFFD33FAD54FFFFFFFFBFFFDFDCCF6F03FFF9FFFFFFFFF45555703967FFFF),
    .INIT_03(256'hFFFFFFF3BEAD5C7FFFFFFFFFFFD794F364B3FFD577FFFFFFF0D55572E167FFFF),
    .INIT_04(256'hFFFFFFF6EC8D551FFFFFFFFFFFF5D751F3E7FFD557FFFFFFF2D555FBC1675FFF),
    .INIT_05(256'hFFFFFFF4EE4D5547FFFFFFFFFFD5D5755EE7FFF57FFFFFFFF15555DBC1673F55),
    .INIT_06(256'hFFFFFFFEDACD5551FFFFFFFFFF5555555F7FFFFD67FFFFFFC3555563CB4506A5),
    .INIT_07(256'hFFFFFFFF30C55556FFFFFFFFF5555555555FFFFDEFFFFFFF6D55554BE347CFD5),
    .INIT_08(256'hFFFFFFFF3C775557A7FFFFFFF5555555555FFFFE1FFFFFFFFD575E6CEBE75BFF),
    .INIT_09(256'hFFFFFFFFC41B5555D27FFF5B75555555557FFFFD7FFFFFFF35555E2CE797DBFF),
    .INIT_0A(256'hFFFFFFFFE61B55555F035DDD55555555555FFFFFFFFFFFFDF55556AF8F37FCFF),
    .INIT_0B(256'hFFFFFFFFF3D3555557DFF555555555555553FFFFFFFFFFFCD5557C2DBD3B75BF),
    .INIT_0C(256'hFFFFFFFFFFD355555555555555555555555CFFFFFFFFFFF7D555720FBC125D3F),
    .INIT_0D(256'hFFFFFFFFFE715555555555555555555555573FFFFFFFFFD355555A8E96D7ED6F),
    .INIT_0E(256'hFFFFFFFFFFF155555555555555555F555555CFFFFFFFFFC75555EA2CF1FEDB6F),
    .INIT_0F(256'hFFFFFFFFFF3B55555555555555557355555573FFFFFFFF6D5555E233CDF67EF3),
    .INIT_10(256'hFFFFFFFFFFA6D555555555555555F3D555555C7FFFFFFD355557C8CF27FF3F3B),
    .INIT_11(256'hFFFFFFFFF6E2D555555555555555F3D555555707FFFFD0D555578FDC9FFF5F46),
    .INIT_12(256'hFFFFFFFFDB70D5555555555555557355555555F8575D0F555557B3705FFFE7F3),
    .INIT_13(256'hFFFFFFFF949455555555555555557D555555557608037D5555548DC1FFFF77F6),
    .INIT_14(256'hFFFFFFDA03165555555555555555555555555557D57D55555555B7AB7FFFD5FE),
    .INIT_15(256'hFFFFFF69DF34F55555555555555557FFF55FD5555555555555555CB217FFFEFF),
    .INIT_16(256'hFFFFFFFFFD3535555555555555FF578000809F5555555555555572FC41FFF57F),
    .INIT_17(256'hFFFFFFFFFCD43555555555FF5C0A82975FFD61D5555555555555CBFD7E2F5F3F),
    .INIT_18(256'hFFFFFFFF526B95555555F582827DFFFFFFFFF6B555555555574763FFFFF67DEF),
    .INIT_19(256'hFFFFFFFEB91F7D555557C09DFFFFFFFFFFFFFF4D55555555572F19FFFFFF5A8B),
    .INIT_1A(256'hFFFFFF8BD8F7CD55555717FFFFFFFFFFFFFFFF735555555555BEDCFFFFFFFD7F),
    .INIT_1B(256'h5555805FD1D5CD55555737FFFFFFFFFFFFFFFF76D55555555E3956FFFFFFFFFF),
    .INIT_1C(256'h559577D55775EF5555579FDDAAA97F7F557DFF7E355555555EAD49BFFFFFFFFF),
    .INIT_1D(256'hFFFFD5557555F35555570A2000000000000AA7722D5555557475689FFFFFFFFF),
    .INIT_1E(256'h555555555557F1D5555708AAAAAAAAAAAAAA8B62875555557051732FFFFFFFFF),
    .INIT_1F(256'h555555555557F8D555572AAAA80022AA0002A2AA835555557E90364FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1125,addra[14:13]}),
    .dia({open_n1129,open_n1130,open_n1131,open_n1132,open_n1133,open_n1134,open_n1135,1'b0,open_n1136}),
    .rsta(rsta),
    .doa({open_n1151,open_n1152,open_n1153,open_n1154,open_n1155,open_n1156,open_n1157,open_n1158,inst_doa_i2_002}));
  // address_offset=16384;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFF7AB8040FFFFFFFB01FFC58444E495EFFCF3FFFFFFF845541318DC0000),
    .INIT_01(256'hFFFFFFCEAAE14AFFFFFFFA0EFFFFBF74BA64BFD8BEFFFFFFF8C554404DCC0000),
    .INIT_02(256'hFFFFFFEBBB6556FFFFFFFCA7FFE6CB7D45FCFFD8F3FFFFFFF405541774395555),
    .INIT_03(256'hFFFFFFEAEB61527FFFFFFFBFFFE2836877FFFFC0B6FFFFFFF955541DA46D1555),
    .INIT_04(256'hFFFFFFF7AFB154BFFFFFFFFFFFC4C70D3EF7FFC117FFFFFFF6155487B12DE100),
    .INIT_05(256'hFFFFFFFEE935152FFFFFFFFFFF05D5404FBFFFD123FFFFFFD5455483A43994FF),
    .INIT_06(256'hFFFFFFFFF965554EFFFFFFFFFC1514555E4FFFD87FFFFFFFFC55547FE13FE6F1),
    .INIT_07(256'hFFFFFFFDAC3555473FFFFFFF90555555512FFFFCAFFFFFFF8155507EC97C7AEA),
    .INIT_08(256'hFFFFFFFFBD345555EBFFFFFCE5555555553FFFF7BFFFFFFFB054530AD9BCDBFF),
    .INIT_09(256'hFFFFFFFF70C855514AAFFFDA55555555550EBFFABFFFFFFFC554539A808C39FF),
    .INIT_0A(256'hFFFFFFFFF748555157EB15C4555555555557BFFFFFFFFFFD8545477AE5C803BF),
    .INIT_0B(256'hFFFFFFFFEDCC5555541FB00555555555555CFFFFFFFFFFFE15454B6AE59DCCBF),
    .INIT_0C(256'hFFFFFFFFF2495550555415545555555555423FFFFFFFFFF315554DAEF2FF73DF),
    .INIT_0D(256'hFFFFFFFFFE195555555555555555515555558EBFFFFFFFED555515BE8431637F),
    .INIT_0E(256'hFFFFFFFFFDDD55555555555555554B55555537BFFFFFFFF1555522BA8D02E8F3),
    .INIT_0F(256'hFFFFFFFFFEDF15555555555555553E15555559FFFFFFFF65555518FA3B5F7B0E),
    .INIT_10(256'hFFFFFFFFFF665555555555555555BA155555433FFFFFFDD55554D6ACFD54EFDD),
    .INIT_11(256'hFFFFFFFFFA8A1555555555555555FA15555554FFFFFFFB5555552A82B0045FF7),
    .INIT_12(256'hFFFFFFFF98CA15555555555555557B15555555327EF5B95555533A1AE4012BCA),
    .INIT_13(256'hFFFFFFFDC70A05555555555555556C5555555542B3EB01555552E82A000583F1),
    .INIT_14(256'hFFFFFFD4ADDF4555555555555550115555555555144015555554F048855473FF),
    .INIT_15(256'hFFFFFFF83F88C55555555555555550001444155555555555555503DCC95406BE),
    .INIT_16(256'hFFFFFFFFFC9C815555555555400443BFFFEED5155555055555554EF228500D3F),
    .INIT_17(256'hFFFFFFFFFA26D155555555004FB13A91FEFA781555555555555427FFB6F1E59F),
    .INIT_18(256'hFFFFFFFFCBFAC555555455AC2B12AFFFFFFFFBD55555555555310EFFFFD7126B),
    .INIT_19(256'hFFFFFFE68CCB25555555AB92FFFFFFFFFFFFFF345555555555F099FFFFFE9ABB),
    .INIT_1A(256'hFFFFFCACA72E615555559FFFFFFFFFFFFFFFFFBD555555555406A2BFFFFFFE02),
    .INIT_1B(256'h0550BF3ECEBF21555545DBFFFFFFFFFFFFFFFFC71555555552D9DE7FFFFFFFFF),
    .INIT_1C(256'h00C15ABFFFFF2C555541D2F5AFAC11904016FFD1855555555133F5FFFFFFFFFF),
    .INIT_1D(256'hAAAABFFFEFFF5955555496D00555500005502F8831555555469FFA6FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFC59555545C11015555555401411B4415555555FE589BFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFF857155545805107EBDD14BFED51C5485555557AAED12FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1184,addra[14:13]}),
    .dia({open_n1188,open_n1189,open_n1190,open_n1191,open_n1192,open_n1193,open_n1194,1'b0,open_n1195}),
    .rsta(rsta),
    .doa({open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,open_n1215,open_n1216,open_n1217,inst_doa_i2_003}));
  // address_offset=16384;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFC8003BE7FFFFFFFCFFFFE75BEE5A793BF7BAFFFFFFFC7FFEE8C36FFFFF),
    .INIT_01(256'hFFFFFFE1000BE5FFFFFFFCF2FFF054DA15C4FFE3FEFFFFFFFC2FFEBF072FFFFF),
    .INIT_02(256'hFFFFFFE5104BF9BFFFFFFE5FFFFD21C3CB56FFE2BEFFFFFFFCEFFEBC57DEAAAA),
    .INIT_03(256'hFFFFFFF5410BF9FFFFFFFFFFFFEC3DC29D57FFEFAFFFFFFFF4FFFEE113DEEAAA),
    .INIT_04(256'hFFFFFFFC011BFE3FFFFFFFFFFFFF3CF2951BFFEEFFFFFFFFE4BFFE21039EFEFF),
    .INIT_05(256'hFFFFFFFD01CFBF9FFFFFFFFFFFBF7FEEF00FFFEEDFFFFFFFE6EFFF74128B7BFF),
    .INIT_06(256'hFFFFFFFD459BFFE7FFFFFFFFFEFFFFFFF1FFFFE7CFFFFFFFC6FFFE80069F095A),
    .INIT_07(256'hFFFFFFFF10CFFFE9FFFFFFFFEFFFFFFFFBFFFFF65BFFFFFFCFFFFA8012DF9BBF),
    .INIT_08(256'hFFFFFFFF14DAFFFF0FFFFFFB0BFFFFFFFFEFFFFC3FFFFFFF1AFFF880060FE3FF),
    .INIT_09(256'hFFFFFFFF9976FFFBF4BFFFF0BFFFFFFFFFEFFFFEFFFFFFFE3FFFFD101A2FF2FF),
    .INIT_0A(256'hFFFFFFFFDD72FFFBFC04AF7EFFFFFFFFFFEFFFFFFFFFFFFE2FFFEC405F2BFDBF),
    .INIT_0B(256'hFFFFFFFFE736FFFFFEA40BAFFFFFFFFFFFE2FFFFFFFFFFF9FFFFE4504F62FE7F),
    .INIT_0C(256'hFFFFFFFFFDB7FFFFFFFEBFFFFFFFFFFFFFEDBFFFFFFFFFFDBFFFE0404971BF7F),
    .INIT_0D(256'hFFFFFFFFFCF6FFFFFFFFFFFFFFFFFEFFFFFF6FFFFFFFFFF3FFFFA4402CFA9FCF),
    .INIT_0E(256'hFFFFFFFFFF67FFFFFFFFFFFFFFFFF5FFFFFFCFFFFFFFFFCFFFFF941077FCF68F),
    .INIT_0F(256'hFFFFFFFFFF30BFFFFFFFFFFFFFFFC5BFFFFFF2FFFFFFFF8FFFFFC54183ADF8B7),
    .INIT_10(256'hFFFFFFFFFE09BFFFFFFFFFFFFFFF44BFFFFFEDFFFFFFFF3FFFFE54064EAB6E66),
    .INIT_11(256'hFFFFFFFFFC10BFFFFFFFFFFFFFFF05BFFFFFFF1BFFFFE5FFFFFF50293FFBAFCC),
    .INIT_12(256'hFFFFFFFFF7A0BFFFFFFFFFFFFFFF85BFFFFFFF90EEEA43FFFFF841E5FBFEDBE0),
    .INIT_13(256'hFFFFFFFE2968EFFFFFFFFFFFFFFFC3FFFFFFFFED1545ABFFFFF90282FFFAEFFD),
    .INIT_14(256'hFFFFFFB0476CEFFFFFFFFFFFFFFFFFFFFFFFFFFFBFEABFFFFFFF4A56BAABBAFC),
    .INIT_15(256'hFFFFFFD2BE3E6FFFFFFFFFFFFFFFFAAABFBEBFFFFFFFFFFFFFFEA9217BABF9FF),
    .INIT_16(256'hFFFFFFFFFF3E6FFFFFFFFFFFEAAFAC4400513FFFFFFFFFFFFFFFE1F9D7FFFEBF),
    .INIT_17(256'hFFFFFFFFF8AD3FFFFFFFFFABB454046BBBFAC7BFFFFFFFFFFFFF87FEBD5BFB3F),
    .INIT_18(256'hFFFFFFFFF1866FFFFFFFFA5411EBBFFFFFFFFD7FFFFFFFFFFF9BD2FFFFB9BECB),
    .INIT_19(256'hFFFFFFFD377ACFFFFFFF003FBFFFFFFFFFFFFFCEFFFFFFFFFF0B76FFFFFFB443),
    .INIT_1A(256'hFFFFFB53B5EE9BFFFFFF7BFFFFFFFFFFFFFFFF83FFFFFFFFFE3C29FFFFFFFEAF),
    .INIT_1B(256'hFFFF51EAA3BFDFFFFFEF6BFFFFFFFFFFFFFFFFF9BFFFFFFFF832ECBFFFFFFFFF),
    .INIT_1C(256'hAA6AFEBFEFFED6FFFFEB2EEA5056EFBEFFAFBFED6FFFFFFFF81BD27FFFFFFFFF),
    .INIT_1D(256'hAAAABFFFEFFFA7FFFFFE51400555500005504FF00BFFFFFFE8BFD17FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFB2FFFFFF040540000000154017D11BFFFFFFF4FEB71FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFA0BFFFFF0504454155540004401006FFFFFFC4646D8BFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1243,addra[14:13]}),
    .dia({open_n1247,open_n1248,open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,1'b0,open_n1254}),
    .rsta(rsta),
    .doa({open_n1269,open_n1270,open_n1271,open_n1272,open_n1273,open_n1274,open_n1275,open_n1276,inst_doa_i2_004}));
  // address_offset=16384;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFDFDDD6BBDFFFDFF68BFFFB0E038C4627CF75FFFFFFF5AAA92CBD2FFFFF),
    .INIT_01(256'hFFFFFFCBFF76B9DFFFFFF22ADFE3D80BD9451FD975FFFFFFF0D2A92820CFFFFF),
    .INIT_02(256'hFFFFFFE7C78E80F57FFFFF8B7FD16F2CC513FDE977FFFFFFF0D2AB8E667FFFFF),
    .INIT_03(256'hFFFFFFDF948CA7B7FFFFDF8D7FFACB1B9281FFE067FFFFFFFB82A95BE4DFFFFF),
    .INIT_04(256'hFFFFFFFAFF3608CFFFFFD5FFFF686B26C767FFC807FFFFFFD04AAB58CE95FFFF),
    .INIT_05(256'hFFFFFFF3FEDAE813FFFFFFFFFD48E8960FA3FFC0237FFFFFF0BAA8A955928D7F),
    .INIT_06(256'hFFFFFFFF199AAA8CFFFFFFFDF7AA2AA88F27FDD82FFFFFFFC52AAA97752D037A),
    .INIT_07(256'hFFFFFFFFD924AA1BFDFFFFFFECAAA2AA8ABFFDC1AFFFFFFF02AAA78945ED4F48),
    .INIT_08(256'hFFFFFFFF4BC7AA80ABFFFFFF30AAAAAAAA9FFFF29FFFFFFF0DA8A627E9D7CFFF),
    .INIT_09(256'hFFFFFFFF2B53AA8E9C1FFFA12AAAAAAAAA3DFF5CB7FFFFFD68AAA1E74BAFD7FF),
    .INIT_0A(256'hFFFFFFFFF9D3AAAE8154DF33AAAAAAAAAA177F57F7FFFFFD728A9F45B0DBFEFF),
    .INIT_0B(256'hFFFFFFFFF0D5AAAAA3EDF25AAAAAAAAAAAA4DF55FFFFFFFDA2AAB0A5913F7CF7),
    .INIT_0C(256'hFFFFFFFFF4E40AAAA0A3C2AAAAAAAAAAAA93B7FFFFFFFFF268AAB58DB7113FBF),
    .INIT_0D(256'hFFFFFFFFFE8EAAAAAAAAAAAAAAAAA0AAAAA06DFFFFFFFFC6AAAAE6AF6E73DF9F),
    .INIT_0E(256'hFFFFFFFFFD3D2AAAAAAAAAAAAAAA8FAAAAAABFFFFFFFFF5CAAAA44456A756F1F),
    .INIT_0F(256'hFFFFFFFFFD43EAAAAAAAAAAAAAAA91EAAAA88DFFFFFFFF88AAAA23F751FD3F71),
    .INIT_10(256'hFFFFFFFFDF4E6AAAAAAAAAAAAAAAF1EAAAA8923FFFFDFC6AAAA3A6D777FFBD1F),
    .INIT_11(256'hFFFFFFF57B3E6AAAAAAAAAAAAAAA7BEAAAAAA0CBFFFFCDAAAAA8BF6F5FF72F83),
    .INIT_12(256'hFFFFFFDF4719CAAAAAAAAAAAAAA8BB6AAAAAAA49898EFEAAAAA71F945FFF77C2),
    .INIT_13(256'hFFFFFDF5E0C93AAAAAAAAAAAAAAAA6AAAAAAAA32C0349EAAAAA7BBFAFFFF5B7B),
    .INIT_14(256'hFFFFFD4D818DDAAAAAAAAAAAAAAAA2AA2AAAAA0AC8BFEAAAAAA38D37BFFF70DF),
    .INIT_15(256'hFFFFFF9C4F9E1AAAAAAAAAAAAA8A275D608BCAAA2A8AAAAAAAA894FB81FF7F7D),
    .INIT_16(256'hFFFFFFFFFE567AAAAAAAAA829F582F2D5DFF1A2AAAAAAAAAAAAA95FA82D5FCB7),
    .INIT_17(256'hFFFFFF7FF4EC62AAAAAAA8D498EAA1CF05DE3DEAAAAAAAAAA80A6FFF7F35F75D),
    .INIT_18(256'hFFFFFFFF201742AAAAA829908D10FFFFFFFFF3C2AAAAAAAAA8BE73FFFF5BAEFF),
    .INIT_19(256'hFFFFFFF7562D18AAAAAA75247FFFFFFFFFFFFF31AAAAAAAAA8C62CFFFFFDA7E7),
    .INIT_1A(256'hFFFFF5E7E471FCAAAAAA4BFFFFFFFFFFFFFFFFC42AAAAAAAA22006FFFFFFFC57),
    .INIT_1B(256'hA2884A2DC24262AAAA9AF3FFFFFFFFFFFFFFFF99EAAAAAAAA650EDFFFFFFDFFF),
    .INIT_1C(256'hA8EA9BE02A00F1AAAAB6A7C4F7D6B595AAFCFFB5FAAAAAAAA6BF545FFFFFFFFF),
    .INIT_1D(256'hFF7F60023003F4AAAAA9EB155AAA2F7FF8A7F31DCC2AAAAAB5BFF46FFFFD7FFF),
    .INIT_1E(256'h0000000000017DAAAAA875557D75F7FF555DEF3550AAAAAAA45E33BFFFFFFFFF),
    .INIT_1F(256'h000000000003DD4AAAA855D762BE00817570755D772AAAAA3A60312F7FFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1302,addra[14:13]}),
    .dia({open_n1306,open_n1307,open_n1308,open_n1309,open_n1310,open_n1311,open_n1312,1'b0,open_n1313}),
    .rsta(rsta),
    .doa({open_n1328,open_n1329,open_n1330,open_n1331,open_n1332,open_n1333,open_n1334,open_n1335,inst_doa_i2_005}));
  // address_offset=16384;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFF08AED74FFFFFFF1F5FFE491DFAFE2FFD1F9FFFFFFF41555EAE7A80000),
    .INIT_01(256'hFFFFFFCAA8C579FFFFFFFDD7FFDAB0EFBB8AFFE7F3FFFFFFF4D5554A55280000),
    .INIT_02(256'hFFFFFFD4804577FFFFFFFC53FFFE11613A54FFCF7BFFFFFFF8B5554D83B80000),
    .INIT_03(256'hFFFFFFF682C555BFFFFFFFFFFFD5B5C95387FFED15FFFFFFF4D557AE21B80000),
    .INIT_04(256'hFFFFFFF02315557FFFFFFFFFFF773E77C623FFCF77FFFFFFD855578C0950A000),
    .INIT_05(256'hFFFFFFFDA19D57FFFFFFFFFFFFD5177BD24FFFEFDBFFFFFFC155572613764AAA),
    .INIT_06(256'hFFFFFFFD087555F7FFFFFFFFFF55555F525FFFC7DBFFFFFFFD55573C915A59F2),
    .INIT_07(256'hFFFFFFFE42E3557FBFFFFFFF595555555D5FFFF757FFFFFF7D555C90979835F7),
    .INIT_08(256'hFFFFFFFFE283555F07FFFFFE2755555555FFFFF3EFFFFFFF2D57561A13B087FF),
    .INIT_09(256'hFFFFFFFF7CE95555EE5FFF4275555555557FFFFDFFFFFFFF75555DDA35080EFF),
    .INIT_0A(256'hFFFFFFFFD92155557CDC080F5555555555C3FFFFFFFFFFFCB57571001DE4037F),
    .INIT_0B(256'hFFFFFFFFDFA5555557F227F555555555557FFFFFFFFFFFFD555573208ECE0A7F),
    .INIT_0C(256'hFFFFFFFFF0DF5555555FFD5555555555557DFFFFFFFFFFF85555766085CFA2EF),
    .INIT_0D(256'hFFFFFFFFFC7F55555555555555555755555F7FFFFFFFFFDF555573A2932292BF),
    .INIT_0E(256'hFFFFFFFFFC36D5555555555555555855555573FFFFFFFFDB555568E23E81D4F3),
    .INIT_0F(256'hFFFFFFFFFD7AD555555555555555EAD5555576FFFFFFFF0D5555DCCA700BB707),
    .INIT_10(256'hFFFFFFFFFFA8555555555555555580D555557FBFFFFFFCF555572A21F000DFEE),
    .INIT_11(256'hFFFFFFFFF52E55555555555555558AD555555F5FFFFFF5D55555F03540022FF3),
    .INIT_12(256'hFFFFFFFF6CC5555555555555555748D555555547BDF87B55555E6AF5200097DC),
    .INIT_13(256'hFFFFFFFECB2F55555555555555557355555555767F545D55555F2555000083F2),
    .INIT_14(256'hFFFFFFE85EC1B5555555555555555D5555555557F57F555555549DE4600023FF),
    .INIT_15(256'hFFFFFFF43F6A1555555555555555DF5D7DDFF555555555555557F5ECEC00097D),
    .INIT_16(256'hFFFFFFFFFC405555555555557F5F52A7FDDF87555555555555555DF514880A3F),
    .INIT_17(256'hFFFFFFFFF717F555555557D7E0F7D568FFF59E555555555555F563FD7BD2824F),
    .INIT_18(256'hFFFFFFFFC7F57D555555FE9FFF255FFFFFFFF5DD55555555577F2DFFFFE92197),
    .INIT_19(256'hFFFFFFDB4CE7AD555557B581FFFFFFFFFFFFFF9F555555555547ECFFFFFD6577),
    .INIT_1A(256'hFFFFFC7E7B1D1555555767FFFFFFFFFFFFFFFFCDD55555555FF4397FFFFFF501),
    .INIT_1B(256'h0AA07F354D7D3D555557C7FFFFFFFFFFFFFFFFC355555555544AA3BFFFFFFFFF),
    .INIT_1C(256'h00C2A57FDFFF3955555701F0FFDC02E02AA9FFE05555555557D22AFFFFFFFFFF),
    .INIT_1D(256'h55557FFDFFFE855555554FCAAAAAAA2AAAA01F4CA5555555736A959FFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFCAED55555622A828A0800AAA02252AF5555557DAE4E7FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFF68B5555554AA83FFFFF7FF57D82C2A5555555E2FDEA9FFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1361,addra[14:13]}),
    .dia({open_n1365,open_n1366,open_n1367,open_n1368,open_n1369,open_n1370,open_n1371,1'b0,open_n1372}),
    .rsta(rsta),
    .doa({open_n1387,open_n1388,open_n1389,open_n1390,open_n1391,open_n1392,open_n1393,open_n1394,inst_doa_i2_006}));
  // address_offset=16384;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFCDDD3FF3FFFFFFF6A2FFF3CFDFF53E17D0F7FFFFFFFCBFFFDFE95FFFFF),
    .INIT_01(256'hFFFFFFDDFD97FEFFFFFFFCA9FFFD67F74CD8FFF8F5FFFFFFFC9FFFF52BDFFFFF),
    .INIT_02(256'hFFFFFFD3D537FC7FFFFFFF8FFFDD745D6789FFDAFDFFFFFFFCFFFF5819EFFFFF),
    .INIT_03(256'hFFFFFFF1D7B7F4FFFFFFFFDFFFFFDCD5ECDBFFF25BFFFFFFF8FFFFD073EFFFFF),
    .INIT_04(256'hFFFFFFFF76C7FFBFFFFFFFFFFFFD5DD9D177FFD28BFFFFFFFB7FFF597B67FFFF),
    .INIT_05(256'hFFFFFFFC74EFFF4FFFFFFFFFFF7FFFFFF7FFFFD287FFFFFFDBFFFF51434797FF),
    .INIT_06(256'hFFFFFFFE5EEFFFD1FFFFFFFFFDFFFFFFF5DFFFD2A7FFFFFFC1FFFD49696F86A5),
    .INIT_07(256'hFFFFFFFFBED7FFF47FFFFFFFDFFFFFFFFFDFFFD22FFFFFFFEFFFFF4D49EFE77F),
    .INIT_08(256'hFFFFFFFF96DFFFFFFFFFFFF55FFFFFFFFF7FFFFC9FFFFFFF5FFFF7676D47F3FF),
    .INIT_09(256'hFFFFFFFF443DFFFFFB7FFFFDFFFFFFFFFFDFFFFFFFFFFFFD3FFFFE8765DFD1FF),
    .INIT_0A(256'hFFFFFFFFE63DFFFFFFA1D57FFFFFFFFFFFFFFFFFFFFFFFFD7FFFF4B5ED97FE7F),
    .INIT_0B(256'hFFFFFFFFD971FFFFFFDD55FFFFFFFFFFFFDBFFFFFFFFFFF4FFFFF4B5DD317DBF),
    .INIT_0C(256'hFFFFFFFFFD7BFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFF57FFFF015D4927FBF),
    .INIT_0D(256'hFFFFFFFFFFF9FFFFFFFFFFFFFFFFFDFFFFFF3FFFFFFFFFFBFFFFDAD7D6F56FCF),
    .INIT_0E(256'hFFFFFFFFFF53FFFFFFFFFFFFFFFFF7FFFFFFEFFFFFFFFFCFFFFF7337F3FCF94F),
    .INIT_0F(256'hFFFFFFFFFF1DFFFFFFFFFFFFFFFF5DFFFFFFF9FFFFFFFF7FFFFFE09D65FEF473),
    .INIT_10(256'hFFFFFFFFFD3F7FFFFFFFFFFFFFFF5DFFFFFFFC7FFFFFFFBFFFFF417D07FF9D99),
    .INIT_11(256'hFFFFFFFFFC497FFFFFFFFFFFFFFF55FFFFFFFFA7FFFFD0FFFFFDA5741FFFDFC4),
    .INIT_12(256'hFFFFFFFFFB527FFFFFFFFFFFFFFF57FFFFFFFF5ADDD527FFFFFD1D527FFFE7D1),
    .INIT_13(256'hFFFFFFFD1696FFFFFFFFFFFFFFFFF5FFFFFFFFFF80A15FFFFFFEFF61FFFFDFFE),
    .INIT_14(256'hFFFFFF708BB4FFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFDD097FFFF5FC),
    .INIT_15(256'hFFFFFFE17D3F5FFFFFFFFFFFFFFFFF5D7F7FFFFFFFFFFFFFFFFDF612B5FFF6FF),
    .INIT_16(256'hFFFFFFFFFF151FFFFFFFFFFFFF5FDDD2A80AD7FFFFFFFFFFFFFFDAF6EBDFFD7F),
    .INIT_17(256'hFFFFFFFFF452BFFFFFFFFFD77782889F77F5CB7FFFFFFFFFFFFF5BFD7CA7FF1F),
    .INIT_18(256'hFFFFFFFFF2499FFFFFFFF7C28AD77FFFFFFFFE1FFFFFFFFFFF6F41FFFF767DC7),
    .INIT_19(256'hFFFFFFFC3B955FFFFFFF48FF7FFFFFFFFFFFFF6FFFFFFFFFFDB73BFFFFFF7883),
    .INIT_1A(256'hFFFFF7815ADD47FFFFFF17FFFFFFFFFFFFFFFFD9FFFFFFFFFDB756FFFFFFFD5F),
    .INIT_1B(256'hFFFFA2D5537FCFFFFFFF17FFFFFFFFFFFFFFFFF47FFFFFFFF73DD47FFFFFFFFF),
    .INIT_1C(256'h5595FD7FDFFDC5FFFFFFDDD50029DFFDD5DF7FDE1FFFFFFFF6A761BFFFFFFFFF),
    .INIT_1D(256'h55557FFFFFFF51FFFFFD288AAAAAAA2AAAA08FF8B7FFFFFFFE7FE2BFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFF7BFFFFFD22000000000000002BE007FFFFFFF0F97B2FFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFD727FFFFD80000AAAAAAAA02A002021FFFFFFD7989E47FFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_016384_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1420,addra[14:13]}),
    .dia({open_n1424,open_n1425,open_n1426,open_n1427,open_n1428,open_n1429,open_n1430,1'b0,open_n1431}),
    .rsta(rsta),
    .doa({open_n1446,open_n1447,open_n1448,open_n1449,open_n1450,open_n1451,open_n1452,open_n1453,inst_doa_i2_007}));
  // address_offset=24576;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hAAAAAAAAAAABFB057DFD1FD78000A020AA80BDDFD7DFFF5FED1545D7FFFFFFFF),
    .INIT_01(256'hAAAAAAAAAAAF531D7DFD7F542AAAAAAAAAAA8B7FFBBFFF5DD7D959737FFFFFFF),
    .INIT_02(256'hAAAAAAAAAA8555197DFFFF5AAAAAAAAAAAAAA83F54BFFF5C9552EE4DFFFFFFFF),
    .INIT_03(256'hAAAAAAAAAAAFEDE05FDD7DC2AAAAAAAAAAAAAA25DF7FFF5815F2AA6813FFFFFF),
    .INIT_04(256'hAAAAAAAAAABF9D73DFDEFDB54AAAAAAAAAAAA8E1DE8FFD59F5F82AAA361FFFFF),
    .INIT_05(256'hAAAAAAAAAA955572B7DEF757E6AAAAAAAAAB1F33564FFF4B55692AAAACE1FFFF),
    .INIT_06(256'hAAAAAAAAAAB6155F4556F6DFF2AAAAAAAAAEFF48FD05FEA955560AAAAAE6DFFF),
    .INIT_07(256'hAAAAAAAAAA77BD572955BCF7F76AAAAAAAABFFF2F68DF2CD55588AAAAA8C79C7),
    .INIT_08(256'hAAAAAAAAAAFEF555CA71DFFFFDA9AAAABA97FFF17215EB0D5572AAAAAAAA792B),
    .INIT_09(256'hAAAAAAAAAAFE555DC31896FFFF74A0008F7FFFFB75FD246D55F4EAAAAAAAA9D2),
    .INIT_0A(256'hAAAAAAAAAA567D5DABCDD87FFFF5FFFF57FFFF555DCEA9E757D6EAAAAAAAAAAB),
    .INIT_0B(256'hAAAAAAAAAA52D55F275DBCFFFFFFFFFFFFFFFF6DDC72276D555A6AAAAAAAAAAA),
    .INIT_0C(256'hAAAAAAAAA877D55F85BFD63FFFFFFFFFFFFFFD5DDECB3F6D555F0AAAAAAAAAAA),
    .INIT_0D(256'hAAAAAAAAA8525557CFF0FAAD7FFFFFFFFFFF5707F73CFF6F5574DAAAAAAAAAAA),
    .INIT_0E(256'hAAAAAAAAA07955574FF303F8757FFFF55D7FDCD5D0B3FFE7557B1AAAAAAAAAAA),
    .INIT_0F(256'hAAAAAAAAA26BD55FCFFA90A102555557F82AD507DDC7FFCF5554BAAAAAAAAAAA),
    .INIT_10(256'hAAAAAAAAAAFF555F8FF774FC357EFF57D55EBB39468FFFCF55CC3AAAAAAAAAAA),
    .INIT_11(256'hAAAAAAAAA809555F0FFC02BF69AAA827C505FDFE2CAFFF4355657AAAAAAAAAAA),
    .INIT_12(256'hAAAAAAAAAA055557AFFE369FFFD5FFFFFFFFFFFE7E3FFF4357887AAAAAAAAAAA),
    .INIT_13(256'hAAAAAAAAA8DD55572FFF155BFFFFFFFFFFFFFFE13EBFFF4B5FA0DAAAAAAAAAAA),
    .INIT_14(256'hAAAAAAAAA90B555F2FFF17C5FFFFFFFFFFFFFD74D8FFFF4354AAEAAAAAAAAAAA),
    .INIT_15(256'hAAAAAAAAAB51D55D2FFF7FF10FFFFFFFFFFFD540F27FFF4B72A86AAAAAAAAAAA),
    .INIT_16(256'hAAAAAAAAA848755D2FFFEBFDE2FF60374227A131EBFFFF67DAA80AAAAAAAAAAA),
    .INIT_17(256'hAAAAAAAAAA5A3D55DFFFC3D828C80AA5F559B887E1FFFF67CAA90AAAAAAAAAAA),
    .INIT_18(256'hAAAAAAAAA5FAAD55DFFFDB7C4BC8020002AB369F2FFFFF4D2AA9AAAAAAAAAAAA),
    .INIT_19(256'hAAAAAAAAAC9AA75DDFFFF9F4ACF71FFD84A2535F0FFFFFC2AAA96AAAAAAAAAAA),
    .INIT_1A(256'hAAAAAAAAA56AA9FD5FFFF9D72987A002662D907C3FFFFFC5AAA9EAAAAAAAAAAA),
    .INIT_1B(256'hAAAAAAAAA0AAAABD5FFFFC976800A1017A55AD5FBFFFFFE1AAA8EAAAAAAAAAAA),
    .INIT_1C(256'h02002A22AF0000A7DFFFFC3DC9A2ADF720578CF8FFFFFF72AAA8580A20800000),
    .INIT_1D(256'h0820002825A88828DFFFFD5D545000A05405A97EFFFFFDFAAAA8902A00002200),
    .INIT_1E(256'h808200A80482820ADFFFFF3DC255005574847FC3FFFFFCE6AAA9500200880222),
    .INIT_1F(256'hAA22AAAA9A682AA6DFFFFF8D71000000000295D3FFFFF2E4AAA9A68A8A2288A8),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1479,addra[14:13]}),
    .dia({open_n1483,open_n1484,open_n1485,open_n1486,open_n1487,open_n1488,open_n1489,1'b0,open_n1490}),
    .rsta(rsta),
    .doa({open_n1505,open_n1506,open_n1507,open_n1508,open_n1509,open_n1510,open_n1511,open_n1512,inst_doa_i3_000}));
  // address_offset=24576;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF4B71AAAA8C0007FFF5FDF557F608002AAAAAA9ACCBD17FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFF882CAAAA8800BD555555555557600096AAAA8FAF3DA597FFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFA2816AAAA00255555555555555740016AAAAA6A8377566FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFD2FAB1AAAA003755555555555555D0002AAAA1AA97FF7DF1FFFFFF),
    .INIT_04(256'hFFFFFFFFFFE2DA86AAA880755555555555555F14029AAA858AB9FFFF533FFFFF),
    .INIT_05(256'hFFFFFFFFFFEA0AA96AA880D7F15555555554FF4E02DAAA0CAA80FFFFF7D9FFFF),
    .INIT_06(256'hFFFFFFFFFF4A6AAB7AA281DFFD5555555553FF57205AAA34AA8ADFFFFF5D67FF),
    .INIT_07(256'hFFFFFFFFFF0BE2AAE6A181F7FC1555555557FFFD82DAA0C8AAA75FFFFFD71F3F),
    .INIT_08(256'hFFFFFFFFFF8BEAAA218789FFFFD4555545F7FFFECB4AA3A8AAAEFFFFFFFF5E3F),
    .INIT_09(256'hFFFFFFFFFF892AA22A6D81FFFF7DFFFFD77FFFF60AEA8E28AA247FFFFFFFFD56),
    .INIT_0A(256'hFFFFFFFFFFA182A2AA9BC57FFFF5FFFF57FFFF7B80D0102AA8277FFFFFFFFFFD),
    .INIT_0B(256'hFFFFFFFFFFA3AAA2AA03DBFFFFFFFFFFFFFFFF78024040A2AAA97FFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFA7AAA22A8B017FFFFFFFFFFFFFFDC602E080A2AAA2DFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFAEAAAAE0298D7D7FFFFFFFFFFF57D023BA00A2AA839FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFF786AAAAE00814A5F57FFFF55D7FF7980B48002AAA8D1FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFF58E2AA2600BF86675FFFFFD557D02502ED0002AAAA41FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFD9EAAA2E00095F6EA010002AAA9DC748AA0002AAA141FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFD7AAAA2E002117FD95557F5E277FDFD116000A6AAB6DFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFAAAAA60026A6FFFFFFFFFFFFFFFFE8A8000A6A85DDFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFD9AAAAA60008A83FFFFFFFFFFFFFFF2290000A6A2F7DFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFDA4AAA26000908B7FFFFFFFFFFFFF37AA0000AEABFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFDE62AA26000080DDFFFFFFFFFFFF9E6AC8000AE87FD7FFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFD7F8AA26000022579802AA0957ABD1CA00000862FFD3FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFD5FC2AA8000262986B5555FF556D0329A00008E3FFDBFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF4DFD2AA8000088B439A0000001F945A800000AE7FFD9FFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF49FF0A28000038A4E419FFD255851AA60000021FFFD1FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF53FFC0280000AAAC92C4AA8F9059BEA80000021FFFD1FFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFDFFFF42800002AAD00A77DC90558EAA80000025FFFD1FFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFF97FFFD8000002E211A00F5D8057A0A20000008FFFFD0FFFDF7FFFFF),
    .INIT_1D(256'hF7DFFFFFF8D777FD000000221C500000540514AA000002AFFFFD8FDDFFFFDDFF),
    .INIT_1E(256'hFFFFFFFFDCFFFFFF000000BAA45500557404428800000197FFFD4FFDFF77FFFF),
    .INIT_1F(256'hFF77FFFFDD7D7FF72000009AAD0000000000D2A00000053DFFFDD7DFDF77DDFD),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1538,addra[14:13]}),
    .dia({open_n1542,open_n1543,open_n1544,open_n1545,open_n1546,open_n1547,open_n1548,1'b0,open_n1549}),
    .rsta(rsta),
    .doa({open_n1564,open_n1565,open_n1566,open_n1567,open_n1568,open_n1569,open_n1570,open_n1571,inst_doa_i3_001}));
  // address_offset=24576;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h555555555557E2755557AAAA0000000000002A2AA9555555471BCAEBFFFFFFFF),
    .INIT_01(256'h55555555555FC7355557AAA800000000000002AAA2D555572FA6F6B6FFFFFFFF),
    .INIT_02(256'h55555555555FED6D5555AAA0000000000000002AA8D555573FC4DD1FBFFFFFFF),
    .INIT_03(256'h55555555555F8FC75555AA88000000000000000AAAD555547FE055D767FFFFFF),
    .INIT_04(256'h55555555557F0FF155552A208000000000000002A8F55552FFE05555FCFFFFFF),
    .INIT_05(256'h55555555557F3FF4D5552A828000000000002A82A835557BFFD255555D87FFFF),
    .INIT_06(256'h55555555557D3FFEB55F288AA00000000000AA208A3557E1FFF8755555D8BFFF),
    .INIT_07(256'h55555555557E3FFF3D5E2AA2A8000000000AAAA0A8B55709FFF07555557DE2DF),
    .INIT_08(256'h5555555555FCBFFFC75C2AAAAA0000000022AAA2B4357C09FFF155555555F742),
    .INIT_09(256'h5555555555FCFFFFC1D422AAAA2A00002A2AAAA2FF15F089FFF9D555555557F5),
    .INIT_0A(256'h5555555555FCFFFF4074222AAAA0AAAA02AAAA2AFF37C28BFFF0D55555555557),
    .INIT_0B(256'h5555555555F4FFFF48BCE8AAAAAAAAAAAAAAAA0BFD9F0A8BFFF4D55555555555),
    .INIT_0C(256'h5555555555FAFFFF4A24F0AAAAAAAAAAAAAAA88BFF3E2A8BFFFE755555555555),
    .INIT_0D(256'h5555555555F1FFFF8A80F0082AAAAAAAAAAA020FDCC0AA8BFFF4F55555555555),
    .INIT_0E(256'h555555555DF3FFFF8AA25AA2A02AAAA0082AA8AFF422AA8BFFF6F55555555555),
    .INIT_0F(256'h555555555DD3FFFF8AA025520AAAAAAAAA80021FF28AAA8BFFFD755555555555),
    .INIT_10(256'h5555555555EBFFFF0AAAE9FD2A000002AAA82277D94AAA8BFFDF755555555555),
    .INIT_11(256'h555555555747FFFF0AA8547FD600000A9F5FFFFD4D0AAA83FFDFB55555555555),
    .INIT_12(256'h55555555554FFFFF0AA83D3FFFFFFFFFFFFFFFFDBD2AAA83FF75B55555555555),
    .INIT_13(256'h5555555557EFFFFF0AAA3FC7FFFFFFFFFFFFFFD67C2AAA83FF5DB55555555555),
    .INIT_14(256'h555555555757FFFF0AAA27DAFFFFFFFFFFFFFFC8F4AAAA83FD55955555555555),
    .INIT_15(256'h5555555557BFFFFF0AAAAFF21FFFFFFFFFFFFE31F0AAAA83F557155555555555),
    .INIT_16(256'h555555555795FFFF0AAA87FAA5FFD55FD57DC2C1D2AAAA8BF557555555555555),
    .INIT_17(256'h5555555555B57FFFAAAA83F4F08000000AA0AFEFC2AAAA8BD557555555555555),
    .INIT_18(256'h555555555FB55FFFAAAAA3FCBC0FFFFFFFC8EB2F4AAAAA8B5557555555555555),
    .INIT_19(256'h555555555D7557FFAAAAA2FD33AAE002F88FAEBF0AAAAA855557D55555555555),
    .INIT_1A(256'h555555555E5555FFAAAAA2FF36F23FFF28FA6EBD2AAAAA8F5557D55555555555),
    .INIT_1B(256'h555555555655557FAAAAA87F8FFF200A8FAA72FE2AAAAA875557D55555555555),
    .INIT_1C(256'h555555555ED5555FAAAAA83FCE5FF002FFA879F4AAAAAAA55557D55555555555),
    .INIT_1D(256'h555555555F555555AAAAAABF63AFFFFFABFAC1F8AAAAAAA55557555555555555),
    .INIT_1E(256'h555555557B555555AAAAAA2FD3AAFFAA8BFBAFD2AAAAA88D5557155555555555),
    .INIT_1F(256'h55DD555571D7D55DAAAAAA0FF2FFFFFFFFFF87EAAAAAA08F55571D7575DD7757),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1597,addra[14:13]}),
    .dia({open_n1601,open_n1602,open_n1603,open_n1604,open_n1605,open_n1606,open_n1607,1'b0,open_n1608}),
    .rsta(rsta),
    .doa({open_n1623,open_n1624,open_n1625,open_n1626,open_n1627,open_n1628,open_n1629,open_n1630,inst_doa_i3_002}));
  // address_offset=24576;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF92A4555450110AFFFFFFFFFFED5115555555560E83E7FFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFF534D555555156FFEAAFFFFFEBF80152155554E4B2A0A3BFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFE416655555155BEFFFFFFFFFFFABC453555542C423FE6CDFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFF4F5644454156BFFFFFFFFFFFFFFF155555547047BFFBEA3FFFFFF),
    .INIT_04(256'hFFFFFFFFFFD5D019055155F0FFFFFFFFFFFFFAFC5585550B5476BFFFE36FFFFF),
    .INIT_05(256'hFFFFFFFFFF80C057555115C3AFFFFFFFFFFFEFF9148554311514BFFFFAF6FFFF),
    .INIT_06(256'hFFFFFFFFFFD18016C152128BFBFFFFFFFFFEFF2E1485569B4001AFFFFFEBCFFF),
    .INIT_07(256'hFFFFFFFFFF93D505B15317B7EBFFFFFFFFFEBFBE514552C6000EEFFFFFFE3E6B),
    .INIT_08(256'hFFFFFFFFFF57D000415313BFFAFFFFFFFEE3FFBC92D52A570119FFFFFFFFBC3F),
    .INIT_09(256'hFFFFFFFFFF12000000164FBFFE3BBAAAEF2FFEBD01C5FD524158FFFFFFFFFEE8),
    .INIT_0A(256'hFFFFFFFFFF02150011068A3FFFE0AFFF03BFFE2241C3A4414147FFFFFFFFFFFE),
    .INIT_0B(256'hFFFFFFFFFE035400455632BFFFFFFFABFAFFFE2000CEC0510007BFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFE1B400145561BEBFFFFFFFFFAFFACAD07B950550005AFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFE4D000185420FF83FFFFFFFFFFE07A406F05514401A6FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFF0C40058551381FE42AAAA0082BFA7517C05551015B2FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFF1D4005C557F59CBAAFFFFABEBBBCF418A1554104487FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFF3D0005C5513AFCC1FFFFF85052F8BD54055545406C3FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFA40005855426FFE2FFFEBBD5FAFEEE63D555494138BFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFA04001D55595CFFFEAFFFFFFFFFFFC0055550915FEBFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFE61000195550073FFFFFFFFFFFFFBE15755550D45FEEFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFE0D000595552947BFFFFFFFFFFEFE3E0515554952FFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFF8840049555155BBFFFFFFFFFFFE6AD1D55555D1BFE7FFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFEAE14049555555A960151007A85BFBF145555594FFF2FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFAF950045554942BC7ABEAFEBAC6A90705555596FFE3FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF8FFF40045555512BE6FAFEFEBF3AAF41555554CBFFE7FFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFC6FF94445555640FBD6AAAEAA7AAA1185555543FFFE3FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFABFFE5405555444BAA8BAAB92FAA8D415555542FFFE7FFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFBFFFFD405555454EAAB8EA17BEAB8455555555AFFFE7FFFFFFFFFFF),
    .INIT_1C(256'hAAAAAFAAF7AAAAF1455554947AAAABFBAAAEA4445555555BFFFE2EAFBAEAAAAA),
    .INIT_1D(256'hAEBAAABEB4FEEEBE45555500FAAAAAFAAAAABF455555555FFFFE2ABFBAAABFAA),
    .INIT_1E(256'hAAAAAAEEB9EAABAF455554351BAAAAAAAAEA94015555567BFFFE7AABAAEEBBAB),
    .INIT_1F(256'hFFFFFFFFEBBFBFFB455555640FAAAAAAAAAA4C0555555B7FFFFEFBFFFFFFFFFE),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1656,addra[14:13]}),
    .dia({open_n1660,open_n1661,open_n1662,open_n1663,open_n1664,open_n1665,open_n1666,1'b0,open_n1667}),
    .rsta(rsta),
    .doa({open_n1682,open_n1683,open_n1684,open_n1685,open_n1686,open_n1687,open_n1688,open_n1689,inst_doa_i3_003}));
  // address_offset=24576;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFAD0AFFFFF4404155555555555140406FFFFFF9F36C083FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFEDF3FFFFF0401554005555541555401BFFFFF4F4DED3CBFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFB9B8BFFFE0005455555555555015101FFFFE87BC9BBEB3FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFEB5ECAEFFE4054555555555555554401BFFFEDFBC1FFBEDAFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFB7FE6AFFB000F5555555555555055002FFFA4EBD4FFFFE9FFFFFF),
    .INIT_05(256'hFFFFFFFFFFFF6FBCFFFB007C5555555555550055406FFE96EAE0FFFFFB4AFFFF),
    .INIT_06(256'hFFFFFFFFFFAF3FEC6FF8057401555555555500D5002FFC17BFE5EFFFFFA43BFF),
    .INIT_07(256'hFFFFFFFFFFAD7AFB1BF804481155555555554045116FF856FFF1AFFFFFFB85BF),
    .INIT_08(256'hFFFFFFFFFFED7FFF8EF9054004155555540C00453C7F8017FEF7FFFFFFFFAF95),
    .INIT_09(256'hFFFFFFFFFFECBFFF92BC514001C1400014D00140FF7F4517BEB2BFFFFFFFFEAB),
    .INIT_0A(256'hFFFFFFFFFFF8EAFFD0AD15C0001F5000FC4001C4FE6C1417BEBDBFFFFFFFFFFE),
    .INIT_0B(256'hFFFFFFFFFFF9EBFF912D904000000054050001C7FE305017FFFCBFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFF1FFFF905DE1140000000005005307FC004013FFF9EFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFB3FFFF1001B047C00000000001FC0BFD440053BFE9EFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFEE3BFFB5004A4551FD5555FF7D4005EF8150017FEACAFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFEE7BFFB10055EE5450000001541416BF4000017FBBAAFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFEC7FFFB5000C2FA15000000550411BAE7D00017BFAAAFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF9FFFFB5001A9BFF95554053BBBFEFF9B500013BEFB6FFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFDFBFFF10013F3FFFFFFFFFFFFFFFFE3F000053EABE6FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFECEFFFF10006F9FFFFFFFFFFFFFFFEDBC000053BBFF6FFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFEFAFFFB10004AE5FFFFFFFFFFFFFFD4FC000017AFFF7FFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFE7BBFFB10000EA12FFFFFFFFFFFFC07F0000007EBFEFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFE3FEBFB10000BB45EBEABAFEFEE0513F0000003BFFFBFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFE2FEAFF400013B8100001554001500BC5000007BFFEEFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFA6FEBFF400006EC404000000040000FC0000017BFFEEFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFAEFFABB400001FF004500000550012F1000001AFFFEAFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF8BFFEAB400005FB100450011540017F4000001AFFFEAFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFDFFFFAB400001FB50014144504000FD4000001AFFFEAFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFCBFFFEE0000017B90000451000006F90000000FFFFEAFFFEFBFFFFF),
    .INIT_1D(256'hFBEFFFFFFAEBBBFE0000003FC0000000000003B50000005FFFFEEFEEEFFFEAFF),
    .INIT_1E(256'hFFFFFFFFF7FFFFFF0000015EF000000000405BE40000004BFFFEFFFEFFBBEFFF),
    .INIT_1F(256'hFFFFFFFFE6BFBFFB1000004FF500000000006FD40000001BFFFE6BFFFFFFFFFE),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1715,addra[14:13]}),
    .dia({open_n1719,open_n1720,open_n1721,open_n1722,open_n1723,open_n1724,open_n1725,1'b0,open_n1726}),
    .rsta(rsta),
    .doa({open_n1741,open_n1742,open_n1743,open_n1744,open_n1745,open_n1746,open_n1747,open_n1748,inst_doa_i3_004}));
  // address_offset=24576;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000029D052AAA815D655FFF5FFFFDD65755C2AAAAABF3DEDD5DFFFFFFF),
    .INIT_01(256'h00000000000DF74A2AA83551554005555541D6D57E6AAA88E57BDBD975FFFFFF),
    .INIT_02(256'h00000000000F5DAEAAAA35CD47DD7FFF55FD0115562AAA1795E8CEE77F7FFFFF),
    .INIT_03(256'h000000000027C7DD1AA255785F5557FD555D5575F70AAA9C3F7882431BFFFFFF),
    .INIT_04(256'h00000000001DBFD05AA7577517555555555758F17F5AAA4D7F7A8002B6BFFFFF),
    .INIT_05(256'h00000000009DD7F922A55E9DED55555555579D3457DAA9017FCB20008C49FFFF),
    .INIT_06(256'h0000000002941FF6D2AF577D59FD55555D5C55E5BDF8A26BFF563000026EDFFF),
    .INIT_07(256'h00000000009D1FFDECACDC7557DF55555559557F3C1A8BEEFF78B0000026F16F),
    .INIT_08(256'h0000000000FEFFFD572578D55717555576BD57F6B3A84CCFFFD800000000712B),
    .INIT_09(256'h0000000000FE7FFDC4613ED555FC0AA8A3D557FEDD6A7EEDFFF66000000021DA),
    .INIT_0A(256'h00000000025657FD0F1BD6D5555557FF755557527F5BF3C7FFDC60000000000B),
    .INIT_0B(256'h0000000002F07FFFA4413CDD555D555555555769D5AF0FCFFFD8400000000000),
    .INIT_0C(256'h0000000000D57FFF0F97DD355555555555555D7D5E14BF47FFF5B00000000000),
    .INIT_0D(256'h000000000AFA7FFF8D7E1DEF5555555555557F1D752DFFCDFFFAD00000000000),
    .INIT_0E(256'h000000000AF1FFFDCD7B0E0E75F5555FF75F761D577355E5FFD9D00000000000),
    .INIT_0F(256'h000000000861FFFD4D58923A6AFD5555482BD605FCA555EFFFD4300000000000),
    .INIT_10(256'h0000000008F5FFFD0D5DD6FFEAFDFFFFAA015D316C0F55EDFF4F300000000000),
    .INIT_11(256'h000000000201FFFDAF5C0A3FE5A003578F87F5DCAD4D55C1FF65D00000000000),
    .INIT_12(256'h0000000002A7FFF50F5E1CBDFF7FD57FFFFFFFFF961555EBFD2A700000000000),
    .INIT_13(256'h00000000035FFFF5AF5DBDFBFFFFFFFFFFFFFFF194B555C3FF08500000000000),
    .INIT_14(256'h000000000321FFFD2F573BED75FFF7FFFFDFFF5DD2D555EBFC20400000000000),
    .INIT_15(256'h00000000035D7FFF25575FF76FFFFFFFFFFFFCBAD8D555EBD023E00000000000),
    .INIT_16(256'h0000000003605FFF255569DC809DF655EA073E57C35D55E5780A800000000000),
    .INIT_17(256'h0000000000729FF7DD55E9DD45B5757F6A050D4549D555CD6801A80000000000),
    .INIT_18(256'h000000000770AFF7FD55F17796D7F7D557347DF7255555EF2001000000000000),
    .INIT_19(256'h000000000C9009FD75557B76DDA4FFFFD93FF6952D5555600801C20200000000),
    .INIT_1A(256'h0000000005A0027DF5557B7D4754C554093F76FE1555554F0801420200000000),
    .INIT_1B(256'h000000000200023D7555543775565DF09FBF52F7355555410803480020880000),
    .INIT_1C(256'h2202AA2A87C8AA8FF55556BDE755D27AD5FF7CF0D55557FA0003680A02000000),
    .INIT_1D(256'h802AA208AD00882275555755F9F555F5FD5F73F6D55557D00003A80A228AAA80),
    .INIT_1E(256'h80AAA028A68A820AF55557B767FF55FFFD1D37C375555CE40001FA202080A2A2),
    .INIT_1F(256'hAAA8AAA81842E824DF5FFD0F7855555555550DFBFD7FF2EEAAA9042220882A8B),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1774,addra[14:13]}),
    .dia({open_n1778,open_n1779,open_n1780,open_n1781,open_n1782,open_n1783,open_n1784,1'b0,open_n1785}),
    .rsta(rsta),
    .doa({open_n1800,open_n1801,open_n1802,open_n1803,open_n1804,open_n1805,open_n1806,open_n1807,inst_doa_i3_005}));
  // address_offset=24576;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF63E1555574AA37F555F555557F80AA9D55555F06C3DBFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFF224F55557CA87D540055555417D2AAA5555574AFB50537FFFFFFF),
    .INIT_02(256'hFFFFFFFFFFDA2A2555574A15455555555555036AA355555CC0B375DCEFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFD8FA31555DAA9055555555555555DAAA75557B0A97FF7F53FFFFFF),
    .INIT_04(256'hFFFFFFFFFFEA72ADD55E28E21555555555555AD6AA9555DDAA917FFDD39FFFFF),
    .INIT_05(256'hFFFFFFFFFF488283555E23880D5555555557A0BF2A55574E2A207FFF75F9FFFF),
    .INIT_06(256'hFFFFFFFFFFE24AAAF55C212801555555555C0007C8555FBEAA027FFFFFD7CFFF),
    .INIT_07(256'hFFFFFFFFFFE3EAAA455CA2200BD5555555580025C2D57CEBAA2DFFFFFFFD3D97),
    .INIT_08(256'hFFFFFFFFFF21CAA8A955040000175555748002AF03F5F2AAAAAEFFFFFFFF5C17),
    .INIT_09(256'hFFFFFFFFFF212AA80B578E0000222002820002A782D50422AA84DFFFFFFFDD54),
    .INIT_0A(256'hFFFFFFFFFD012AA8A8554400000002AA00000224A8DE30A0AA8FDFFFFFFFFFFD),
    .INIT_0B(256'hFFFFFFFFFD83AAA8809D7608000800000000020EA230C2A8AA837FFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFDA7AAA88A890D8000000000000008BEA0A32A28AAAA7FFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFF8E2AA88A8BC5480000000000000290A322AAAAAAAF9FFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFF8CAAAA4AA21D56A0000000000A82F28BE2AA82AAA79FFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFF2EAAAACAABF8E76202AAA00A89FFF88792AA82AA849FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFF3EAAAACAA21DFCDDFDFFF5FFDFF676828AAA8AAA961FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF58AAAA4AA813FF7BDFFF778055FDFD302AAA86AA14FFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFF2AAA2EAAA62EFFFD57FFFFFFFFFFEC82AAAA6AAFD5FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFF92AAA26AAA00ABFFFFFFFFFFFFFFFA2BAAAA8EA8FDDFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFD2EAAAA6AAA1E037FFFFFFFFFFFFDBF0A2AAAAEA9DFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFD4CAAA86AAA22AFDFFFFFFFFFFFD0AE2EAAAAA6A7DFDFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFF7D2AA86AAAAAACBBCA28889FD83EBC28AAAAA687F71FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFF5FEAA08AAA86898EF55FF5E00CE090B0AAAAAEBFFDBFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF4DFD2A08AAA8A2B0A320000021CAA582AAAAAAC7FFDBFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF49FFEA88AAAA9A26A9AAAAA2B70A2624AAAAAA3F7FD3DFDFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF5FFFFA80AAAA8A842254AA8BF0A29422AAAAA81F7FDBDFDFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFF7FFFFE80AAAA8807808F5D5D0AA092AAAAAAAA5F7FFBFFFDF77FFFF),
    .INIT_1C(256'h5555555579DD55728AAAA8683A00005A00AA0808AAAAA88FFFFF355577D55555),
    .INIT_1D(256'hDD7FD775D8FDDD5D8AAAA80018A00000A80A9E8AAAAAAAAFFFFF357777DFFFD5),
    .INIT_1E(256'h555555D5F6DD555F8AAAAABA04AA00AAA808A802AAAAA917FFFDEF7775DD75D5),
    .INIT_1F(256'hFFFFFFFFD77FFFF78AAAAA9A060000000002E80AAAAAA59FFFFDF7FFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1833,addra[14:13]}),
    .dia({open_n1837,open_n1838,open_n1839,open_n1840,open_n1841,open_n1842,open_n1843,1'b0,open_n1844}),
    .rsta(rsta),
    .doa({open_n1859,open_n1860,open_n1861,open_n1862,open_n1863,open_n1864,open_n1865,open_n1866,inst_doa_i3_006}));
  // address_offset=24576;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFF5E3DFFFFF0000000000000000200003FFFFFF67B1C043FFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFDE3BFFFFF800800155000001402000B7FFFFF3F84DE3C7FFFFFFF),
    .INIT_02(256'hFFFFFFFFFFF56757FFFD80201000000000005400007FFFFD3F6677973FFFFFFF),
    .INIT_03(256'hFFFFFFFFFFD7ADEDFFFD000F000000000000000000FFFFFCF5C2FF7FE5FFFFFF),
    .INIT_04(256'hFFFFFFFFFFF7AD53FFFF001F4000000000000580025FFFD8D5E8FFFFD6FFFFFF),
    .INIT_05(256'hFFFFFFFFFFF79D7E7FFF0077F800000000025FE2021FFF51D5D0FFFFF785FFFF),
    .INIT_06(256'hFFFFFFFFFF5F355F1FFD00D7F4000000000BFFF0009FFF4355DAFFFFFF5837FF),
    .INIT_07(256'hFFFFFFFFFFDEB55797FF83DFF6800000000FFFD0A21FFD0B55D27FFFFFF74A7F),
    .INIT_08(256'hFFFFFFFFFFDEB5576DF409FFFDC20000215FFD50FE3FF5AB5573FFFFFFFF5F6A),
    .INIT_09(256'hFFFFFFFFFFDC555769768BFFFFD7D55575FFFD527F3FD22B55717FFFFFFFFD57),
    .INIT_0A(256'hFFFFFFFFFFF4D557E8DC03FFFFFFFD55FFFFFDDBD515682B557A7FFFFFFFFFFD),
    .INIT_0B(256'hFFFFFFFFFF76D557683C49F7FFF7FFFFFFFFFDF95FD52023557C7FFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFF72D55760A4D8FFFFFFFFFFFFFFF7635D5680A35556FFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFD73D557E008F837FFFFFFFFFFFFFD475C520023555CDFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFD535557A00858A35FFFFFFFFFF5558D7E88002B555CDFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFDDB5557200AAD701F5555555FF4A81772C0002B55755FFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFDCB5557A000E1F722A8AAAA0028887DDBE0002B55575FFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFF6F5557A002547FDC0000A0F777FDFF4520002355F71FFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFF4D555F20023F1FFFFFFFFFFFFFFFFFBF800003557D9FFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFCD555F20009F67FFFFFFFFFFFFFFF67C00002357FF9FFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFDD5555720008DDAFFFFFFFFFFFFFF42FC00000357FFBFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFDBF555720000D589FFFFFFFFFFFFF51F000000B57FFBFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFF1FD55720000773CDF57FD7D55D6B4BF00000037FFF7FFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFD1F555F8000237E5AAAAAA01FF83547CA0000035FFD5FFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFF59FD55F800009DED50D555555637D8FC000000B7FFDDFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFF5DFFD57800002DD9DE37FFF5E25F79F20000005FFFD5FFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFF4FFFF5780000AD7975295554A5F74BD80000025FFFD5FFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFEFFFF57800002FFA55588A285FF56DE80000025FFFF5FFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFCF7FFDD000002B747555D0755FF51F600000007FFFF7FFFDD7FFFFF),
    .INIT_1D(256'h77D57DFF75D777FD0000003FC5F55555FD5F637A000000AFFFFFFFDDDD75557F),
    .INIT_1E(256'hFFFFFFFF7BF7FFFF0000002DF9FF55FFFD5DC7D800000087FFFDB5DDDF77DF7F),
    .INIT_1F(256'hFFFFFFFFD97FFFF72000008DFB55555555553FE800000027FFFD97FFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32768x8_sub_024576_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1892,addra[14:13]}),
    .dia({open_n1896,open_n1897,open_n1898,open_n1899,open_n1900,open_n1901,open_n1902,1'b0,open_n1903}),
    .rsta(rsta),
    .doa({open_n1918,open_n1919,open_n1920,open_n1921,open_n1922,open_n1923,open_n1924,open_n1925,inst_doa_i3_007}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(doa[7]));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

